// This is the unpowered netlist.
module spell (clock,
    i_la_wb_disable,
    i_la_write,
    i_wb_cyc,
    i_wb_stb,
    i_wb_we,
    interrupt,
    o_wb_ack,
    rambus_wb_ack_i,
    rambus_wb_clk_o,
    rambus_wb_cyc_o,
    rambus_wb_rst_o,
    rambus_wb_stb_o,
    rambus_wb_we_o,
    reset,
    i_la_addr,
    i_la_data,
    i_wb_addr,
    i_wb_data,
    io_in,
    io_oeb,
    io_out,
    la_data_out,
    o_wb_data,
    rambus_wb_addr_o,
    rambus_wb_dat_i,
    rambus_wb_dat_o,
    rambus_wb_sel_o);
 input clock;
 input i_la_wb_disable;
 input i_la_write;
 input i_wb_cyc;
 input i_wb_stb;
 input i_wb_we;
 output interrupt;
 output o_wb_ack;
 input rambus_wb_ack_i;
 output rambus_wb_clk_o;
 output rambus_wb_cyc_o;
 output rambus_wb_rst_o;
 output rambus_wb_stb_o;
 output rambus_wb_we_o;
 input reset;
 input [6:0] i_la_addr;
 input [7:0] i_la_data;
 input [31:0] i_wb_addr;
 input [31:0] i_wb_data;
 input [7:0] io_in;
 output [7:0] io_oeb;
 output [7:0] io_out;
 output [31:0] la_data_out;
 output [31:0] o_wb_data;
 output [9:0] rambus_wb_addr_o;
 input [31:0] rambus_wb_dat_i;
 output [31:0] rambus_wb_dat_o;
 output [3:0] rambus_wb_sel_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire \cycles_per_ms[0] ;
 wire \cycles_per_ms[10] ;
 wire \cycles_per_ms[11] ;
 wire \cycles_per_ms[12] ;
 wire \cycles_per_ms[13] ;
 wire \cycles_per_ms[14] ;
 wire \cycles_per_ms[15] ;
 wire \cycles_per_ms[16] ;
 wire \cycles_per_ms[17] ;
 wire \cycles_per_ms[18] ;
 wire \cycles_per_ms[19] ;
 wire \cycles_per_ms[1] ;
 wire \cycles_per_ms[20] ;
 wire \cycles_per_ms[21] ;
 wire \cycles_per_ms[22] ;
 wire \cycles_per_ms[23] ;
 wire \cycles_per_ms[2] ;
 wire \cycles_per_ms[3] ;
 wire \cycles_per_ms[4] ;
 wire \cycles_per_ms[5] ;
 wire \cycles_per_ms[6] ;
 wire \cycles_per_ms[7] ;
 wire \cycles_per_ms[8] ;
 wire \cycles_per_ms[9] ;
 wire \delay_counter[0] ;
 wire \delay_counter[1] ;
 wire \delay_counter[2] ;
 wire \delay_counter[3] ;
 wire \delay_counter[4] ;
 wire \delay_counter[5] ;
 wire \delay_counter[6] ;
 wire \delay_counter[7] ;
 wire \delay_cycles[0] ;
 wire \delay_cycles[10] ;
 wire \delay_cycles[11] ;
 wire \delay_cycles[12] ;
 wire \delay_cycles[13] ;
 wire \delay_cycles[14] ;
 wire \delay_cycles[15] ;
 wire \delay_cycles[16] ;
 wire \delay_cycles[17] ;
 wire \delay_cycles[18] ;
 wire \delay_cycles[19] ;
 wire \delay_cycles[1] ;
 wire \delay_cycles[20] ;
 wire \delay_cycles[21] ;
 wire \delay_cycles[22] ;
 wire \delay_cycles[23] ;
 wire \delay_cycles[2] ;
 wire \delay_cycles[3] ;
 wire \delay_cycles[4] ;
 wire \delay_cycles[5] ;
 wire \delay_cycles[6] ;
 wire \delay_cycles[7] ;
 wire \delay_cycles[8] ;
 wire \delay_cycles[9] ;
 wire edge_interrupts;
 wire \exec.memory_input[0] ;
 wire \exec.memory_input[1] ;
 wire \exec.memory_input[2] ;
 wire \exec.memory_input[3] ;
 wire \exec.memory_input[4] ;
 wire \exec.memory_input[5] ;
 wire \exec.memory_input[6] ;
 wire \exec.memory_input[7] ;
 wire \exec.out_of_order_exec ;
 wire \intr[0] ;
 wire \intr[1] ;
 wire \intr_enable[0] ;
 wire \intr_enable[1] ;
 wire \mem.addr[0] ;
 wire \mem.addr[1] ;
 wire \mem.dff_data_out[0] ;
 wire \mem.dff_data_out[1] ;
 wire \mem.dff_data_out[2] ;
 wire \mem.dff_data_out[3] ;
 wire \mem.dff_data_out[4] ;
 wire \mem.dff_data_out[5] ;
 wire \mem.dff_data_out[6] ;
 wire \mem.dff_data_out[7] ;
 wire \mem.dff_data_ready ;
 wire \mem.io_data_out[0] ;
 wire \mem.io_data_out[1] ;
 wire \mem.io_data_out[2] ;
 wire \mem.io_data_out[3] ;
 wire \mem.io_data_out[4] ;
 wire \mem.io_data_out[5] ;
 wire \mem.io_data_out[6] ;
 wire \mem.io_data_out[7] ;
 wire \mem.io_data_ready ;
 wire \mem.mem_dff.code_mem[0][0] ;
 wire \mem.mem_dff.code_mem[0][1] ;
 wire \mem.mem_dff.code_mem[0][2] ;
 wire \mem.mem_dff.code_mem[0][3] ;
 wire \mem.mem_dff.code_mem[0][4] ;
 wire \mem.mem_dff.code_mem[0][5] ;
 wire \mem.mem_dff.code_mem[0][6] ;
 wire \mem.mem_dff.code_mem[0][7] ;
 wire \mem.mem_dff.code_mem[10][0] ;
 wire \mem.mem_dff.code_mem[10][1] ;
 wire \mem.mem_dff.code_mem[10][2] ;
 wire \mem.mem_dff.code_mem[10][3] ;
 wire \mem.mem_dff.code_mem[10][4] ;
 wire \mem.mem_dff.code_mem[10][5] ;
 wire \mem.mem_dff.code_mem[10][6] ;
 wire \mem.mem_dff.code_mem[10][7] ;
 wire \mem.mem_dff.code_mem[11][0] ;
 wire \mem.mem_dff.code_mem[11][1] ;
 wire \mem.mem_dff.code_mem[11][2] ;
 wire \mem.mem_dff.code_mem[11][3] ;
 wire \mem.mem_dff.code_mem[11][4] ;
 wire \mem.mem_dff.code_mem[11][5] ;
 wire \mem.mem_dff.code_mem[11][6] ;
 wire \mem.mem_dff.code_mem[11][7] ;
 wire \mem.mem_dff.code_mem[12][0] ;
 wire \mem.mem_dff.code_mem[12][1] ;
 wire \mem.mem_dff.code_mem[12][2] ;
 wire \mem.mem_dff.code_mem[12][3] ;
 wire \mem.mem_dff.code_mem[12][4] ;
 wire \mem.mem_dff.code_mem[12][5] ;
 wire \mem.mem_dff.code_mem[12][6] ;
 wire \mem.mem_dff.code_mem[12][7] ;
 wire \mem.mem_dff.code_mem[13][0] ;
 wire \mem.mem_dff.code_mem[13][1] ;
 wire \mem.mem_dff.code_mem[13][2] ;
 wire \mem.mem_dff.code_mem[13][3] ;
 wire \mem.mem_dff.code_mem[13][4] ;
 wire \mem.mem_dff.code_mem[13][5] ;
 wire \mem.mem_dff.code_mem[13][6] ;
 wire \mem.mem_dff.code_mem[13][7] ;
 wire \mem.mem_dff.code_mem[14][0] ;
 wire \mem.mem_dff.code_mem[14][1] ;
 wire \mem.mem_dff.code_mem[14][2] ;
 wire \mem.mem_dff.code_mem[14][3] ;
 wire \mem.mem_dff.code_mem[14][4] ;
 wire \mem.mem_dff.code_mem[14][5] ;
 wire \mem.mem_dff.code_mem[14][6] ;
 wire \mem.mem_dff.code_mem[14][7] ;
 wire \mem.mem_dff.code_mem[15][0] ;
 wire \mem.mem_dff.code_mem[15][1] ;
 wire \mem.mem_dff.code_mem[15][2] ;
 wire \mem.mem_dff.code_mem[15][3] ;
 wire \mem.mem_dff.code_mem[15][4] ;
 wire \mem.mem_dff.code_mem[15][5] ;
 wire \mem.mem_dff.code_mem[15][6] ;
 wire \mem.mem_dff.code_mem[15][7] ;
 wire \mem.mem_dff.code_mem[16][0] ;
 wire \mem.mem_dff.code_mem[16][1] ;
 wire \mem.mem_dff.code_mem[16][2] ;
 wire \mem.mem_dff.code_mem[16][3] ;
 wire \mem.mem_dff.code_mem[16][4] ;
 wire \mem.mem_dff.code_mem[16][5] ;
 wire \mem.mem_dff.code_mem[16][6] ;
 wire \mem.mem_dff.code_mem[16][7] ;
 wire \mem.mem_dff.code_mem[17][0] ;
 wire \mem.mem_dff.code_mem[17][1] ;
 wire \mem.mem_dff.code_mem[17][2] ;
 wire \mem.mem_dff.code_mem[17][3] ;
 wire \mem.mem_dff.code_mem[17][4] ;
 wire \mem.mem_dff.code_mem[17][5] ;
 wire \mem.mem_dff.code_mem[17][6] ;
 wire \mem.mem_dff.code_mem[17][7] ;
 wire \mem.mem_dff.code_mem[18][0] ;
 wire \mem.mem_dff.code_mem[18][1] ;
 wire \mem.mem_dff.code_mem[18][2] ;
 wire \mem.mem_dff.code_mem[18][3] ;
 wire \mem.mem_dff.code_mem[18][4] ;
 wire \mem.mem_dff.code_mem[18][5] ;
 wire \mem.mem_dff.code_mem[18][6] ;
 wire \mem.mem_dff.code_mem[18][7] ;
 wire \mem.mem_dff.code_mem[19][0] ;
 wire \mem.mem_dff.code_mem[19][1] ;
 wire \mem.mem_dff.code_mem[19][2] ;
 wire \mem.mem_dff.code_mem[19][3] ;
 wire \mem.mem_dff.code_mem[19][4] ;
 wire \mem.mem_dff.code_mem[19][5] ;
 wire \mem.mem_dff.code_mem[19][6] ;
 wire \mem.mem_dff.code_mem[19][7] ;
 wire \mem.mem_dff.code_mem[1][0] ;
 wire \mem.mem_dff.code_mem[1][1] ;
 wire \mem.mem_dff.code_mem[1][2] ;
 wire \mem.mem_dff.code_mem[1][3] ;
 wire \mem.mem_dff.code_mem[1][4] ;
 wire \mem.mem_dff.code_mem[1][5] ;
 wire \mem.mem_dff.code_mem[1][6] ;
 wire \mem.mem_dff.code_mem[1][7] ;
 wire \mem.mem_dff.code_mem[20][0] ;
 wire \mem.mem_dff.code_mem[20][1] ;
 wire \mem.mem_dff.code_mem[20][2] ;
 wire \mem.mem_dff.code_mem[20][3] ;
 wire \mem.mem_dff.code_mem[20][4] ;
 wire \mem.mem_dff.code_mem[20][5] ;
 wire \mem.mem_dff.code_mem[20][6] ;
 wire \mem.mem_dff.code_mem[20][7] ;
 wire \mem.mem_dff.code_mem[21][0] ;
 wire \mem.mem_dff.code_mem[21][1] ;
 wire \mem.mem_dff.code_mem[21][2] ;
 wire \mem.mem_dff.code_mem[21][3] ;
 wire \mem.mem_dff.code_mem[21][4] ;
 wire \mem.mem_dff.code_mem[21][5] ;
 wire \mem.mem_dff.code_mem[21][6] ;
 wire \mem.mem_dff.code_mem[21][7] ;
 wire \mem.mem_dff.code_mem[22][0] ;
 wire \mem.mem_dff.code_mem[22][1] ;
 wire \mem.mem_dff.code_mem[22][2] ;
 wire \mem.mem_dff.code_mem[22][3] ;
 wire \mem.mem_dff.code_mem[22][4] ;
 wire \mem.mem_dff.code_mem[22][5] ;
 wire \mem.mem_dff.code_mem[22][6] ;
 wire \mem.mem_dff.code_mem[22][7] ;
 wire \mem.mem_dff.code_mem[23][0] ;
 wire \mem.mem_dff.code_mem[23][1] ;
 wire \mem.mem_dff.code_mem[23][2] ;
 wire \mem.mem_dff.code_mem[23][3] ;
 wire \mem.mem_dff.code_mem[23][4] ;
 wire \mem.mem_dff.code_mem[23][5] ;
 wire \mem.mem_dff.code_mem[23][6] ;
 wire \mem.mem_dff.code_mem[23][7] ;
 wire \mem.mem_dff.code_mem[24][0] ;
 wire \mem.mem_dff.code_mem[24][1] ;
 wire \mem.mem_dff.code_mem[24][2] ;
 wire \mem.mem_dff.code_mem[24][3] ;
 wire \mem.mem_dff.code_mem[24][4] ;
 wire \mem.mem_dff.code_mem[24][5] ;
 wire \mem.mem_dff.code_mem[24][6] ;
 wire \mem.mem_dff.code_mem[24][7] ;
 wire \mem.mem_dff.code_mem[25][0] ;
 wire \mem.mem_dff.code_mem[25][1] ;
 wire \mem.mem_dff.code_mem[25][2] ;
 wire \mem.mem_dff.code_mem[25][3] ;
 wire \mem.mem_dff.code_mem[25][4] ;
 wire \mem.mem_dff.code_mem[25][5] ;
 wire \mem.mem_dff.code_mem[25][6] ;
 wire \mem.mem_dff.code_mem[25][7] ;
 wire \mem.mem_dff.code_mem[26][0] ;
 wire \mem.mem_dff.code_mem[26][1] ;
 wire \mem.mem_dff.code_mem[26][2] ;
 wire \mem.mem_dff.code_mem[26][3] ;
 wire \mem.mem_dff.code_mem[26][4] ;
 wire \mem.mem_dff.code_mem[26][5] ;
 wire \mem.mem_dff.code_mem[26][6] ;
 wire \mem.mem_dff.code_mem[26][7] ;
 wire \mem.mem_dff.code_mem[27][0] ;
 wire \mem.mem_dff.code_mem[27][1] ;
 wire \mem.mem_dff.code_mem[27][2] ;
 wire \mem.mem_dff.code_mem[27][3] ;
 wire \mem.mem_dff.code_mem[27][4] ;
 wire \mem.mem_dff.code_mem[27][5] ;
 wire \mem.mem_dff.code_mem[27][6] ;
 wire \mem.mem_dff.code_mem[27][7] ;
 wire \mem.mem_dff.code_mem[28][0] ;
 wire \mem.mem_dff.code_mem[28][1] ;
 wire \mem.mem_dff.code_mem[28][2] ;
 wire \mem.mem_dff.code_mem[28][3] ;
 wire \mem.mem_dff.code_mem[28][4] ;
 wire \mem.mem_dff.code_mem[28][5] ;
 wire \mem.mem_dff.code_mem[28][6] ;
 wire \mem.mem_dff.code_mem[28][7] ;
 wire \mem.mem_dff.code_mem[29][0] ;
 wire \mem.mem_dff.code_mem[29][1] ;
 wire \mem.mem_dff.code_mem[29][2] ;
 wire \mem.mem_dff.code_mem[29][3] ;
 wire \mem.mem_dff.code_mem[29][4] ;
 wire \mem.mem_dff.code_mem[29][5] ;
 wire \mem.mem_dff.code_mem[29][6] ;
 wire \mem.mem_dff.code_mem[29][7] ;
 wire \mem.mem_dff.code_mem[2][0] ;
 wire \mem.mem_dff.code_mem[2][1] ;
 wire \mem.mem_dff.code_mem[2][2] ;
 wire \mem.mem_dff.code_mem[2][3] ;
 wire \mem.mem_dff.code_mem[2][4] ;
 wire \mem.mem_dff.code_mem[2][5] ;
 wire \mem.mem_dff.code_mem[2][6] ;
 wire \mem.mem_dff.code_mem[2][7] ;
 wire \mem.mem_dff.code_mem[30][0] ;
 wire \mem.mem_dff.code_mem[30][1] ;
 wire \mem.mem_dff.code_mem[30][2] ;
 wire \mem.mem_dff.code_mem[30][3] ;
 wire \mem.mem_dff.code_mem[30][4] ;
 wire \mem.mem_dff.code_mem[30][5] ;
 wire \mem.mem_dff.code_mem[30][6] ;
 wire \mem.mem_dff.code_mem[30][7] ;
 wire \mem.mem_dff.code_mem[31][0] ;
 wire \mem.mem_dff.code_mem[31][1] ;
 wire \mem.mem_dff.code_mem[31][2] ;
 wire \mem.mem_dff.code_mem[31][3] ;
 wire \mem.mem_dff.code_mem[31][4] ;
 wire \mem.mem_dff.code_mem[31][5] ;
 wire \mem.mem_dff.code_mem[31][6] ;
 wire \mem.mem_dff.code_mem[31][7] ;
 wire \mem.mem_dff.code_mem[3][0] ;
 wire \mem.mem_dff.code_mem[3][1] ;
 wire \mem.mem_dff.code_mem[3][2] ;
 wire \mem.mem_dff.code_mem[3][3] ;
 wire \mem.mem_dff.code_mem[3][4] ;
 wire \mem.mem_dff.code_mem[3][5] ;
 wire \mem.mem_dff.code_mem[3][6] ;
 wire \mem.mem_dff.code_mem[3][7] ;
 wire \mem.mem_dff.code_mem[4][0] ;
 wire \mem.mem_dff.code_mem[4][1] ;
 wire \mem.mem_dff.code_mem[4][2] ;
 wire \mem.mem_dff.code_mem[4][3] ;
 wire \mem.mem_dff.code_mem[4][4] ;
 wire \mem.mem_dff.code_mem[4][5] ;
 wire \mem.mem_dff.code_mem[4][6] ;
 wire \mem.mem_dff.code_mem[4][7] ;
 wire \mem.mem_dff.code_mem[5][0] ;
 wire \mem.mem_dff.code_mem[5][1] ;
 wire \mem.mem_dff.code_mem[5][2] ;
 wire \mem.mem_dff.code_mem[5][3] ;
 wire \mem.mem_dff.code_mem[5][4] ;
 wire \mem.mem_dff.code_mem[5][5] ;
 wire \mem.mem_dff.code_mem[5][6] ;
 wire \mem.mem_dff.code_mem[5][7] ;
 wire \mem.mem_dff.code_mem[6][0] ;
 wire \mem.mem_dff.code_mem[6][1] ;
 wire \mem.mem_dff.code_mem[6][2] ;
 wire \mem.mem_dff.code_mem[6][3] ;
 wire \mem.mem_dff.code_mem[6][4] ;
 wire \mem.mem_dff.code_mem[6][5] ;
 wire \mem.mem_dff.code_mem[6][6] ;
 wire \mem.mem_dff.code_mem[6][7] ;
 wire \mem.mem_dff.code_mem[7][0] ;
 wire \mem.mem_dff.code_mem[7][1] ;
 wire \mem.mem_dff.code_mem[7][2] ;
 wire \mem.mem_dff.code_mem[7][3] ;
 wire \mem.mem_dff.code_mem[7][4] ;
 wire \mem.mem_dff.code_mem[7][5] ;
 wire \mem.mem_dff.code_mem[7][6] ;
 wire \mem.mem_dff.code_mem[7][7] ;
 wire \mem.mem_dff.code_mem[8][0] ;
 wire \mem.mem_dff.code_mem[8][1] ;
 wire \mem.mem_dff.code_mem[8][2] ;
 wire \mem.mem_dff.code_mem[8][3] ;
 wire \mem.mem_dff.code_mem[8][4] ;
 wire \mem.mem_dff.code_mem[8][5] ;
 wire \mem.mem_dff.code_mem[8][6] ;
 wire \mem.mem_dff.code_mem[8][7] ;
 wire \mem.mem_dff.code_mem[9][0] ;
 wire \mem.mem_dff.code_mem[9][1] ;
 wire \mem.mem_dff.code_mem[9][2] ;
 wire \mem.mem_dff.code_mem[9][3] ;
 wire \mem.mem_dff.code_mem[9][4] ;
 wire \mem.mem_dff.code_mem[9][5] ;
 wire \mem.mem_dff.code_mem[9][6] ;
 wire \mem.mem_dff.code_mem[9][7] ;
 wire \mem.mem_dff.cycles[0] ;
 wire \mem.mem_dff.cycles[1] ;
 wire \mem.mem_dff.data_mem[0][0] ;
 wire \mem.mem_dff.data_mem[0][1] ;
 wire \mem.mem_dff.data_mem[0][2] ;
 wire \mem.mem_dff.data_mem[0][3] ;
 wire \mem.mem_dff.data_mem[0][4] ;
 wire \mem.mem_dff.data_mem[0][5] ;
 wire \mem.mem_dff.data_mem[0][6] ;
 wire \mem.mem_dff.data_mem[0][7] ;
 wire \mem.mem_dff.data_mem[1][0] ;
 wire \mem.mem_dff.data_mem[1][1] ;
 wire \mem.mem_dff.data_mem[1][2] ;
 wire \mem.mem_dff.data_mem[1][3] ;
 wire \mem.mem_dff.data_mem[1][4] ;
 wire \mem.mem_dff.data_mem[1][5] ;
 wire \mem.mem_dff.data_mem[1][6] ;
 wire \mem.mem_dff.data_mem[1][7] ;
 wire \mem.mem_dff.data_mem[2][0] ;
 wire \mem.mem_dff.data_mem[2][1] ;
 wire \mem.mem_dff.data_mem[2][2] ;
 wire \mem.mem_dff.data_mem[2][3] ;
 wire \mem.mem_dff.data_mem[2][4] ;
 wire \mem.mem_dff.data_mem[2][5] ;
 wire \mem.mem_dff.data_mem[2][6] ;
 wire \mem.mem_dff.data_mem[2][7] ;
 wire \mem.mem_dff.data_mem[3][0] ;
 wire \mem.mem_dff.data_mem[3][1] ;
 wire \mem.mem_dff.data_mem[3][2] ;
 wire \mem.mem_dff.data_mem[3][3] ;
 wire \mem.mem_dff.data_mem[3][4] ;
 wire \mem.mem_dff.data_mem[3][5] ;
 wire \mem.mem_dff.data_mem[3][6] ;
 wire \mem.mem_dff.data_mem[3][7] ;
 wire \mem.mem_dff.data_mem[4][0] ;
 wire \mem.mem_dff.data_mem[4][1] ;
 wire \mem.mem_dff.data_mem[4][2] ;
 wire \mem.mem_dff.data_mem[4][3] ;
 wire \mem.mem_dff.data_mem[4][4] ;
 wire \mem.mem_dff.data_mem[4][5] ;
 wire \mem.mem_dff.data_mem[4][6] ;
 wire \mem.mem_dff.data_mem[4][7] ;
 wire \mem.mem_dff.data_mem[5][0] ;
 wire \mem.mem_dff.data_mem[5][1] ;
 wire \mem.mem_dff.data_mem[5][2] ;
 wire \mem.mem_dff.data_mem[5][3] ;
 wire \mem.mem_dff.data_mem[5][4] ;
 wire \mem.mem_dff.data_mem[5][5] ;
 wire \mem.mem_dff.data_mem[5][6] ;
 wire \mem.mem_dff.data_mem[5][7] ;
 wire \mem.mem_dff.data_mem[6][0] ;
 wire \mem.mem_dff.data_mem[6][1] ;
 wire \mem.mem_dff.data_mem[6][2] ;
 wire \mem.mem_dff.data_mem[6][3] ;
 wire \mem.mem_dff.data_mem[6][4] ;
 wire \mem.mem_dff.data_mem[6][5] ;
 wire \mem.mem_dff.data_mem[6][6] ;
 wire \mem.mem_dff.data_mem[6][7] ;
 wire \mem.mem_dff.data_mem[7][0] ;
 wire \mem.mem_dff.data_mem[7][1] ;
 wire \mem.mem_dff.data_mem[7][2] ;
 wire \mem.mem_dff.data_mem[7][3] ;
 wire \mem.mem_dff.data_mem[7][4] ;
 wire \mem.mem_dff.data_mem[7][5] ;
 wire \mem.mem_dff.data_mem[7][6] ;
 wire \mem.mem_dff.data_mem[7][7] ;
 wire \mem.mem_dff.memory_type_data ;
 wire \mem.mem_io.past_write ;
 wire \mem.select ;
 wire \mem.sram_enable ;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire prev_level_interrupt;
 wire prev_reg_write;
 wire net268;
 wire net269;
 wire clknet_leaf_0_clock;
 wire single_step;
 wire \stack[0][0] ;
 wire \stack[0][1] ;
 wire \stack[0][2] ;
 wire \stack[0][3] ;
 wire \stack[0][4] ;
 wire \stack[0][5] ;
 wire \stack[0][6] ;
 wire \stack[0][7] ;
 wire \stack[10][0] ;
 wire \stack[10][1] ;
 wire \stack[10][2] ;
 wire \stack[10][3] ;
 wire \stack[10][4] ;
 wire \stack[10][5] ;
 wire \stack[10][6] ;
 wire \stack[10][7] ;
 wire \stack[11][0] ;
 wire \stack[11][1] ;
 wire \stack[11][2] ;
 wire \stack[11][3] ;
 wire \stack[11][4] ;
 wire \stack[11][5] ;
 wire \stack[11][6] ;
 wire \stack[11][7] ;
 wire \stack[12][0] ;
 wire \stack[12][1] ;
 wire \stack[12][2] ;
 wire \stack[12][3] ;
 wire \stack[12][4] ;
 wire \stack[12][5] ;
 wire \stack[12][6] ;
 wire \stack[12][7] ;
 wire \stack[13][0] ;
 wire \stack[13][1] ;
 wire \stack[13][2] ;
 wire \stack[13][3] ;
 wire \stack[13][4] ;
 wire \stack[13][5] ;
 wire \stack[13][6] ;
 wire \stack[13][7] ;
 wire \stack[14][0] ;
 wire \stack[14][1] ;
 wire \stack[14][2] ;
 wire \stack[14][3] ;
 wire \stack[14][4] ;
 wire \stack[14][5] ;
 wire \stack[14][6] ;
 wire \stack[14][7] ;
 wire \stack[15][0] ;
 wire \stack[15][1] ;
 wire \stack[15][2] ;
 wire \stack[15][3] ;
 wire \stack[15][4] ;
 wire \stack[15][5] ;
 wire \stack[15][6] ;
 wire \stack[15][7] ;
 wire \stack[16][0] ;
 wire \stack[16][1] ;
 wire \stack[16][2] ;
 wire \stack[16][3] ;
 wire \stack[16][4] ;
 wire \stack[16][5] ;
 wire \stack[16][6] ;
 wire \stack[16][7] ;
 wire \stack[17][0] ;
 wire \stack[17][1] ;
 wire \stack[17][2] ;
 wire \stack[17][3] ;
 wire \stack[17][4] ;
 wire \stack[17][5] ;
 wire \stack[17][6] ;
 wire \stack[17][7] ;
 wire \stack[18][0] ;
 wire \stack[18][1] ;
 wire \stack[18][2] ;
 wire \stack[18][3] ;
 wire \stack[18][4] ;
 wire \stack[18][5] ;
 wire \stack[18][6] ;
 wire \stack[18][7] ;
 wire \stack[19][0] ;
 wire \stack[19][1] ;
 wire \stack[19][2] ;
 wire \stack[19][3] ;
 wire \stack[19][4] ;
 wire \stack[19][5] ;
 wire \stack[19][6] ;
 wire \stack[19][7] ;
 wire \stack[1][0] ;
 wire \stack[1][1] ;
 wire \stack[1][2] ;
 wire \stack[1][3] ;
 wire \stack[1][4] ;
 wire \stack[1][5] ;
 wire \stack[1][6] ;
 wire \stack[1][7] ;
 wire \stack[20][0] ;
 wire \stack[20][1] ;
 wire \stack[20][2] ;
 wire \stack[20][3] ;
 wire \stack[20][4] ;
 wire \stack[20][5] ;
 wire \stack[20][6] ;
 wire \stack[20][7] ;
 wire \stack[21][0] ;
 wire \stack[21][1] ;
 wire \stack[21][2] ;
 wire \stack[21][3] ;
 wire \stack[21][4] ;
 wire \stack[21][5] ;
 wire \stack[21][6] ;
 wire \stack[21][7] ;
 wire \stack[22][0] ;
 wire \stack[22][1] ;
 wire \stack[22][2] ;
 wire \stack[22][3] ;
 wire \stack[22][4] ;
 wire \stack[22][5] ;
 wire \stack[22][6] ;
 wire \stack[22][7] ;
 wire \stack[23][0] ;
 wire \stack[23][1] ;
 wire \stack[23][2] ;
 wire \stack[23][3] ;
 wire \stack[23][4] ;
 wire \stack[23][5] ;
 wire \stack[23][6] ;
 wire \stack[23][7] ;
 wire \stack[24][0] ;
 wire \stack[24][1] ;
 wire \stack[24][2] ;
 wire \stack[24][3] ;
 wire \stack[24][4] ;
 wire \stack[24][5] ;
 wire \stack[24][6] ;
 wire \stack[24][7] ;
 wire \stack[25][0] ;
 wire \stack[25][1] ;
 wire \stack[25][2] ;
 wire \stack[25][3] ;
 wire \stack[25][4] ;
 wire \stack[25][5] ;
 wire \stack[25][6] ;
 wire \stack[25][7] ;
 wire \stack[26][0] ;
 wire \stack[26][1] ;
 wire \stack[26][2] ;
 wire \stack[26][3] ;
 wire \stack[26][4] ;
 wire \stack[26][5] ;
 wire \stack[26][6] ;
 wire \stack[26][7] ;
 wire \stack[27][0] ;
 wire \stack[27][1] ;
 wire \stack[27][2] ;
 wire \stack[27][3] ;
 wire \stack[27][4] ;
 wire \stack[27][5] ;
 wire \stack[27][6] ;
 wire \stack[27][7] ;
 wire \stack[28][0] ;
 wire \stack[28][1] ;
 wire \stack[28][2] ;
 wire \stack[28][3] ;
 wire \stack[28][4] ;
 wire \stack[28][5] ;
 wire \stack[28][6] ;
 wire \stack[28][7] ;
 wire \stack[29][0] ;
 wire \stack[29][1] ;
 wire \stack[29][2] ;
 wire \stack[29][3] ;
 wire \stack[29][4] ;
 wire \stack[29][5] ;
 wire \stack[29][6] ;
 wire \stack[29][7] ;
 wire \stack[2][0] ;
 wire \stack[2][1] ;
 wire \stack[2][2] ;
 wire \stack[2][3] ;
 wire \stack[2][4] ;
 wire \stack[2][5] ;
 wire \stack[2][6] ;
 wire \stack[2][7] ;
 wire \stack[30][0] ;
 wire \stack[30][1] ;
 wire \stack[30][2] ;
 wire \stack[30][3] ;
 wire \stack[30][4] ;
 wire \stack[30][5] ;
 wire \stack[30][6] ;
 wire \stack[30][7] ;
 wire \stack[31][0] ;
 wire \stack[31][1] ;
 wire \stack[31][2] ;
 wire \stack[31][3] ;
 wire \stack[31][4] ;
 wire \stack[31][5] ;
 wire \stack[31][6] ;
 wire \stack[31][7] ;
 wire \stack[3][0] ;
 wire \stack[3][1] ;
 wire \stack[3][2] ;
 wire \stack[3][3] ;
 wire \stack[3][4] ;
 wire \stack[3][5] ;
 wire \stack[3][6] ;
 wire \stack[3][7] ;
 wire \stack[4][0] ;
 wire \stack[4][1] ;
 wire \stack[4][2] ;
 wire \stack[4][3] ;
 wire \stack[4][4] ;
 wire \stack[4][5] ;
 wire \stack[4][6] ;
 wire \stack[4][7] ;
 wire \stack[5][0] ;
 wire \stack[5][1] ;
 wire \stack[5][2] ;
 wire \stack[5][3] ;
 wire \stack[5][4] ;
 wire \stack[5][5] ;
 wire \stack[5][6] ;
 wire \stack[5][7] ;
 wire \stack[6][0] ;
 wire \stack[6][1] ;
 wire \stack[6][2] ;
 wire \stack[6][3] ;
 wire \stack[6][4] ;
 wire \stack[6][5] ;
 wire \stack[6][6] ;
 wire \stack[6][7] ;
 wire \stack[7][0] ;
 wire \stack[7][1] ;
 wire \stack[7][2] ;
 wire \stack[7][3] ;
 wire \stack[7][4] ;
 wire \stack[7][5] ;
 wire \stack[7][6] ;
 wire \stack[7][7] ;
 wire \stack[8][0] ;
 wire \stack[8][1] ;
 wire \stack[8][2] ;
 wire \stack[8][3] ;
 wire \stack[8][4] ;
 wire \stack[8][5] ;
 wire \stack[8][6] ;
 wire \stack[8][7] ;
 wire \stack[9][0] ;
 wire \stack[9][1] ;
 wire \stack[9][2] ;
 wire \stack[9][3] ;
 wire \stack[9][4] ;
 wire \stack[9][5] ;
 wire \stack[9][6] ;
 wire \stack[9][7] ;
 wire wb_read_ack;
 wire wb_write_ack;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire clknet_leaf_3_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_6_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_20_clock;
 wire clknet_leaf_21_clock;
 wire clknet_leaf_22_clock;
 wire clknet_leaf_23_clock;
 wire clknet_leaf_24_clock;
 wire clknet_leaf_25_clock;
 wire clknet_leaf_26_clock;
 wire clknet_leaf_29_clock;
 wire clknet_leaf_30_clock;
 wire clknet_leaf_31_clock;
 wire clknet_leaf_32_clock;
 wire clknet_leaf_33_clock;
 wire clknet_leaf_34_clock;
 wire clknet_leaf_35_clock;
 wire clknet_leaf_36_clock;
 wire clknet_leaf_37_clock;
 wire clknet_leaf_38_clock;
 wire clknet_leaf_39_clock;
 wire clknet_leaf_40_clock;
 wire clknet_leaf_41_clock;
 wire clknet_leaf_42_clock;
 wire clknet_leaf_43_clock;
 wire clknet_leaf_44_clock;
 wire clknet_leaf_45_clock;
 wire clknet_leaf_46_clock;
 wire clknet_leaf_47_clock;
 wire clknet_leaf_48_clock;
 wire clknet_leaf_49_clock;
 wire clknet_leaf_50_clock;
 wire clknet_leaf_51_clock;
 wire clknet_leaf_53_clock;
 wire clknet_leaf_54_clock;
 wire clknet_leaf_55_clock;
 wire clknet_leaf_56_clock;
 wire clknet_leaf_57_clock;
 wire clknet_leaf_58_clock;
 wire clknet_leaf_59_clock;
 wire clknet_leaf_60_clock;
 wire clknet_leaf_61_clock;
 wire clknet_leaf_62_clock;
 wire clknet_leaf_64_clock;
 wire clknet_leaf_65_clock;
 wire clknet_leaf_66_clock;
 wire clknet_leaf_67_clock;
 wire clknet_leaf_68_clock;
 wire clknet_leaf_69_clock;
 wire clknet_leaf_70_clock;
 wire clknet_leaf_71_clock;
 wire clknet_leaf_72_clock;
 wire clknet_leaf_73_clock;
 wire clknet_leaf_74_clock;
 wire clknet_leaf_75_clock;
 wire clknet_leaf_76_clock;
 wire clknet_leaf_77_clock;
 wire clknet_leaf_78_clock;
 wire clknet_leaf_79_clock;
 wire clknet_leaf_80_clock;
 wire clknet_leaf_81_clock;
 wire clknet_leaf_82_clock;
 wire clknet_leaf_84_clock;
 wire clknet_leaf_85_clock;
 wire clknet_leaf_86_clock;
 wire clknet_leaf_87_clock;
 wire clknet_leaf_88_clock;
 wire clknet_leaf_89_clock;
 wire clknet_leaf_90_clock;
 wire clknet_leaf_91_clock;
 wire clknet_leaf_92_clock;
 wire clknet_leaf_93_clock;
 wire clknet_leaf_94_clock;
 wire clknet_leaf_95_clock;
 wire clknet_leaf_96_clock;
 wire clknet_leaf_97_clock;
 wire clknet_leaf_98_clock;
 wire clknet_leaf_99_clock;
 wire clknet_leaf_100_clock;
 wire clknet_leaf_101_clock;
 wire clknet_leaf_102_clock;
 wire clknet_leaf_103_clock;
 wire clknet_leaf_104_clock;
 wire clknet_leaf_105_clock;
 wire clknet_leaf_106_clock;
 wire clknet_leaf_107_clock;
 wire clknet_leaf_108_clock;
 wire clknet_leaf_109_clock;
 wire clknet_leaf_110_clock;
 wire clknet_leaf_111_clock;
 wire clknet_leaf_112_clock;
 wire clknet_leaf_113_clock;
 wire clknet_leaf_114_clock;
 wire clknet_leaf_115_clock;
 wire clknet_leaf_116_clock;
 wire clknet_leaf_117_clock;
 wire clknet_leaf_118_clock;
 wire clknet_leaf_119_clock;
 wire clknet_leaf_120_clock;
 wire clknet_leaf_122_clock;
 wire clknet_leaf_123_clock;
 wire clknet_leaf_124_clock;
 wire clknet_leaf_125_clock;
 wire clknet_leaf_127_clock;
 wire clknet_leaf_128_clock;
 wire clknet_leaf_129_clock;
 wire clknet_leaf_131_clock;
 wire clknet_leaf_132_clock;
 wire clknet_leaf_133_clock;
 wire clknet_leaf_134_clock;
 wire clknet_leaf_135_clock;
 wire clknet_leaf_138_clock;
 wire clknet_leaf_139_clock;
 wire clknet_leaf_140_clock;
 wire clknet_leaf_141_clock;
 wire clknet_leaf_142_clock;
 wire clknet_leaf_143_clock;
 wire clknet_leaf_144_clock;
 wire clknet_leaf_145_clock;
 wire clknet_leaf_146_clock;
 wire clknet_leaf_147_clock;
 wire clknet_leaf_148_clock;
 wire clknet_leaf_149_clock;
 wire clknet_leaf_150_clock;
 wire clknet_leaf_151_clock;
 wire clknet_leaf_152_clock;
 wire clknet_leaf_153_clock;
 wire clknet_leaf_154_clock;
 wire clknet_leaf_156_clock;
 wire clknet_leaf_157_clock;
 wire clknet_leaf_158_clock;
 wire clknet_leaf_159_clock;
 wire clknet_leaf_160_clock;
 wire clknet_leaf_161_clock;
 wire clknet_leaf_162_clock;
 wire clknet_leaf_163_clock;
 wire clknet_leaf_166_clock;
 wire clknet_leaf_167_clock;
 wire clknet_leaf_168_clock;
 wire clknet_leaf_169_clock;
 wire clknet_leaf_170_clock;
 wire clknet_leaf_171_clock;
 wire clknet_leaf_173_clock;
 wire clknet_leaf_175_clock;
 wire clknet_leaf_176_clock;
 wire clknet_leaf_177_clock;
 wire clknet_leaf_178_clock;
 wire clknet_leaf_179_clock;
 wire clknet_leaf_180_clock;
 wire clknet_leaf_181_clock;
 wire clknet_leaf_182_clock;
 wire clknet_leaf_183_clock;
 wire clknet_leaf_184_clock;
 wire clknet_leaf_185_clock;
 wire clknet_leaf_186_clock;
 wire clknet_leaf_187_clock;
 wire clknet_leaf_188_clock;
 wire clknet_leaf_189_clock;
 wire clknet_leaf_190_clock;
 wire clknet_leaf_191_clock;
 wire clknet_leaf_192_clock;
 wire clknet_leaf_193_clock;
 wire clknet_0_clock;
 wire clknet_2_0_0_clock;
 wire clknet_2_1_0_clock;
 wire clknet_2_2_0_clock;
 wire clknet_2_3_0_clock;
 wire clknet_3_0_0_clock;
 wire clknet_3_1_0_clock;
 wire clknet_3_2_0_clock;
 wire clknet_3_3_0_clock;
 wire clknet_3_4_0_clock;
 wire clknet_3_5_0_clock;
 wire clknet_3_6_0_clock;
 wire clknet_3_7_0_clock;
 wire clknet_4_0_0_clock;
 wire clknet_4_1_0_clock;
 wire clknet_4_2_0_clock;
 wire clknet_4_3_0_clock;
 wire clknet_4_4_0_clock;
 wire clknet_4_5_0_clock;
 wire clknet_4_6_0_clock;
 wire clknet_4_7_0_clock;
 wire clknet_4_8_0_clock;
 wire clknet_4_9_0_clock;
 wire clknet_4_10_0_clock;
 wire clknet_4_11_0_clock;
 wire clknet_4_12_0_clock;
 wire clknet_4_13_0_clock;
 wire clknet_4_14_0_clock;
 wire clknet_4_15_0_clock;
 wire clknet_opt_1_0_clock;
 wire clknet_opt_2_0_clock;
 wire clknet_opt_3_0_clock;
 wire clknet_opt_4_0_clock;
 wire clknet_opt_4_1_clock;
 wire clknet_opt_5_0_clock;
 wire clknet_opt_6_0_clock;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05196_ (.I(\mem.addr[1] ),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05197_ (.I(\mem.addr[0] ),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05198_ (.A1(_00756_),
    .A2(_00757_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05199_ (.I(_00758_),
    .ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05200_ (.A1(\mem.addr[1] ),
    .A2(\mem.addr[0] ),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05201_ (.I(_00759_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05202_ (.I(_00760_),
    .ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05203_ (.A1(\mem.addr[1] ),
    .A2(_00757_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05204_ (.I(_00761_),
    .ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05205_ (.A1(_00756_),
    .A2(\mem.addr[0] ),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05206_ (.I(_00762_),
    .ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05207_ (.I(\mem.select ),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05208_ (.I(\mem.mem_dff.memory_type_data ),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05209_ (.A1(_00763_),
    .A2(_00764_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05210_ (.I(_00765_),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05211_ (.I(net136),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05212_ (.I(_00766_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05213_ (.I(net135),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05214_ (.I(_00768_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05215_ (.I(_00769_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05216_ (.A1(_00767_),
    .A2(_00770_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05217_ (.I(_00771_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05218_ (.I(net138),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05219_ (.I(net137),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05220_ (.I(net136),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05221_ (.A1(_00773_),
    .A2(_00774_),
    .A3(_00775_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05222_ (.A1(net140),
    .A2(_00776_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05223_ (.I(net140),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05224_ (.A1(_00778_),
    .A2(_00771_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05225_ (.A1(_00772_),
    .A2(_00777_),
    .B(_00779_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05226_ (.I(_00780_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05227_ (.A1(_00774_),
    .A2(_00775_),
    .A3(_00768_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05228_ (.I(_00782_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05229_ (.I(_00775_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05230_ (.I(net135),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05231_ (.I(net137),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05232_ (.A1(_00784_),
    .A2(_00785_),
    .B(_00786_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05233_ (.A1(_00783_),
    .A2(_00787_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05234_ (.I(_00788_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05235_ (.I(net135),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05236_ (.I(_00790_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05237_ (.I(_00791_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05238_ (.I(_00784_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05239_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05240_ (.I0(\stack[3][0] ),
    .I1(\stack[0][0] ),
    .I2(\stack[1][0] ),
    .I3(\stack[2][0] ),
    .S0(_00792_),
    .S1(_00794_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05241_ (.A1(_00789_),
    .A2(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05242_ (.I(_00787_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05243_ (.A1(_00783_),
    .A2(_00797_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05244_ (.I(_00798_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05245_ (.I(_00769_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05246_ (.I(_00800_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05247_ (.I(_00766_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05248_ (.I(_00802_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05249_ (.I0(\stack[7][0] ),
    .I1(\stack[4][0] ),
    .I2(\stack[5][0] ),
    .I3(\stack[6][0] ),
    .S0(_00801_),
    .S1(_00803_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05250_ (.I(net138),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05251_ (.A1(_00805_),
    .A2(_00782_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05252_ (.I(_00806_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05253_ (.A1(_00799_),
    .A2(_00804_),
    .B(_00807_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05254_ (.I(_00785_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05255_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05256_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05257_ (.I0(\stack[11][0] ),
    .I1(\stack[8][0] ),
    .I2(\stack[9][0] ),
    .I3(\stack[10][0] ),
    .S0(_00811_),
    .S1(_00794_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05258_ (.A1(_00789_),
    .A2(_00812_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05259_ (.I0(\stack[15][0] ),
    .I1(\stack[12][0] ),
    .I2(\stack[13][0] ),
    .I3(\stack[14][0] ),
    .S0(_00801_),
    .S1(_00803_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05260_ (.A1(_00773_),
    .A2(_00782_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05261_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05262_ (.A1(_00799_),
    .A2(_00814_),
    .B(_00816_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05263_ (.A1(_00796_),
    .A2(_00808_),
    .B1(_00813_),
    .B2(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05264_ (.I(_00798_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05265_ (.I(_00768_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05266_ (.I(_00820_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05267_ (.I(_00821_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05268_ (.I(_00802_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05269_ (.I0(\stack[31][0] ),
    .I1(\stack[28][0] ),
    .I2(\stack[29][0] ),
    .I3(\stack[30][0] ),
    .S0(_00822_),
    .S1(_00823_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05270_ (.I(_00783_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05271_ (.I(_00797_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05272_ (.I(_00769_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05273_ (.I(_00784_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05274_ (.I0(\stack[27][0] ),
    .I1(\stack[24][0] ),
    .I2(\stack[25][0] ),
    .I3(\stack[26][0] ),
    .S0(_00827_),
    .S1(_00828_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05275_ (.A1(_00825_),
    .A2(_00826_),
    .A3(_00829_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05276_ (.A1(_00819_),
    .A2(_00824_),
    .B(_00830_),
    .C(_00816_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05277_ (.I(_00827_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05278_ (.I0(\stack[23][0] ),
    .I1(\stack[20][0] ),
    .I2(\stack[21][0] ),
    .I3(\stack[22][0] ),
    .S0(_00832_),
    .S1(_00823_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05279_ (.I0(\stack[19][0] ),
    .I1(\stack[16][0] ),
    .I2(\stack[17][0] ),
    .I3(\stack[18][0] ),
    .S0(_00821_),
    .S1(_00828_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05280_ (.A1(_00825_),
    .A2(_00826_),
    .A3(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05281_ (.A1(_00819_),
    .A2(_00833_),
    .B(_00835_),
    .C(_00807_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05282_ (.A1(_00831_),
    .A2(_00836_),
    .B(_00781_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05283_ (.A1(_00781_),
    .A2(_00818_),
    .B(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05284_ (.I(_00838_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05285_ (.I(_00839_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05286_ (.I(_00840_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05287_ (.I(_00841_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05288_ (.I(_00842_),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05289_ (.I(_00810_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05290_ (.I(_00793_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05291_ (.I0(\stack[19][1] ),
    .I1(\stack[16][1] ),
    .I2(\stack[17][1] ),
    .I3(\stack[18][1] ),
    .S0(_00843_),
    .S1(_00844_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05292_ (.A1(_00789_),
    .A2(_00845_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05293_ (.I(_00802_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05294_ (.I0(\stack[23][1] ),
    .I1(\stack[20][1] ),
    .I2(\stack[21][1] ),
    .I3(\stack[22][1] ),
    .S0(_00822_),
    .S1(_00847_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05295_ (.A1(_00819_),
    .A2(_00848_),
    .B(_00807_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05296_ (.I(net140),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05297_ (.A1(_00850_),
    .A2(_00776_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05298_ (.I(_00851_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05299_ (.A1(_00850_),
    .A2(_00772_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05300_ (.A1(_00772_),
    .A2(_00852_),
    .B(_00853_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05301_ (.I(_00768_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05302_ (.I(_00855_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05303_ (.I(_00856_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05304_ (.I0(\stack[31][1] ),
    .I1(\stack[28][1] ),
    .I2(\stack[29][1] ),
    .I3(\stack[30][1] ),
    .S0(_00857_),
    .S1(_00847_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05305_ (.I0(\stack[27][1] ),
    .I1(\stack[24][1] ),
    .I2(\stack[25][1] ),
    .I3(\stack[26][1] ),
    .S0(_00856_),
    .S1(_00793_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05306_ (.A1(_00783_),
    .A2(_00797_),
    .A3(_00859_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05307_ (.A1(_00798_),
    .A2(_00858_),
    .B(_00860_),
    .C(_00816_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05308_ (.A1(_00846_),
    .A2(_00849_),
    .B(_00854_),
    .C(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05309_ (.I0(\stack[3][1] ),
    .I1(\stack[0][1] ),
    .I2(\stack[1][1] ),
    .I3(\stack[2][1] ),
    .S0(_00811_),
    .S1(_00794_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05310_ (.A1(_00789_),
    .A2(_00863_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05311_ (.I0(\stack[7][1] ),
    .I1(\stack[4][1] ),
    .I2(\stack[5][1] ),
    .I3(\stack[6][1] ),
    .S0(_00832_),
    .S1(_00823_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05312_ (.A1(_00819_),
    .A2(_00865_),
    .B(_00807_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05313_ (.I0(\stack[15][1] ),
    .I1(\stack[12][1] ),
    .I2(\stack[13][1] ),
    .I3(\stack[14][1] ),
    .S0(_00857_),
    .S1(_00847_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05314_ (.I(_00855_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05315_ (.I(_00784_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05316_ (.I0(\stack[11][1] ),
    .I1(\stack[8][1] ),
    .I2(\stack[9][1] ),
    .I3(\stack[10][1] ),
    .S0(_00868_),
    .S1(_00869_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05317_ (.A1(_00825_),
    .A2(_00797_),
    .A3(_00870_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05318_ (.A1(_00798_),
    .A2(_00867_),
    .B(_00871_),
    .C(_00816_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05319_ (.A1(_00864_),
    .A2(_00866_),
    .B(_00780_),
    .C(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05320_ (.A1(_00862_),
    .A2(_00873_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05321_ (.I(_00874_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05322_ (.I(_00875_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05323_ (.I(_00876_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05324_ (.I(_00877_),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05325_ (.I(_00806_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05326_ (.I(_00878_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05327_ (.I(_00785_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05328_ (.I(_00880_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05329_ (.I(_00881_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05330_ (.I(_00767_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05331_ (.I(_00883_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05332_ (.I0(\stack[31][2] ),
    .I1(\stack[28][2] ),
    .I2(\stack[29][2] ),
    .I3(\stack[30][2] ),
    .S0(_00882_),
    .S1(_00884_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05333_ (.I0(\stack[27][2] ),
    .I1(\stack[24][2] ),
    .I2(\stack[25][2] ),
    .I3(\stack[26][2] ),
    .S0(_00882_),
    .S1(_00884_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05334_ (.I(_00788_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05335_ (.I0(_00885_),
    .I1(_00886_),
    .S(_00887_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05336_ (.I(_00887_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05337_ (.I(_00767_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05338_ (.I(_00890_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05339_ (.I0(\stack[19][2] ),
    .I1(\stack[16][2] ),
    .I2(\stack[17][2] ),
    .I3(\stack[18][2] ),
    .S0(_00843_),
    .S1(_00891_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05340_ (.I(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05341_ (.I(_00825_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05342_ (.I0(\stack[23][2] ),
    .I1(\stack[20][2] ),
    .I2(\stack[21][2] ),
    .I3(\stack[22][2] ),
    .S0(_00822_),
    .S1(_00823_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05343_ (.A1(_00894_),
    .A2(_00826_),
    .B(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05344_ (.A1(_00889_),
    .A2(_00893_),
    .B(_00896_),
    .C(_00878_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05345_ (.A1(_00879_),
    .A2(_00888_),
    .B(_00897_),
    .C(_00854_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05346_ (.I(_00785_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05347_ (.I(_00899_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05348_ (.I(_00900_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05349_ (.I(_00883_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05350_ (.I0(\stack[11][2] ),
    .I1(\stack[8][2] ),
    .I2(\stack[9][2] ),
    .I3(\stack[10][2] ),
    .S0(_00901_),
    .S1(_00902_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05351_ (.I(_00903_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05352_ (.I(_00826_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05353_ (.I0(\stack[15][2] ),
    .I1(\stack[12][2] ),
    .I2(\stack[13][2] ),
    .I3(\stack[14][2] ),
    .S0(_00843_),
    .S1(_00891_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05354_ (.A1(_00894_),
    .A2(_00905_),
    .B(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05355_ (.I(_00815_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05356_ (.A1(_00889_),
    .A2(_00904_),
    .B(_00907_),
    .C(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05357_ (.I0(\stack[3][2] ),
    .I1(\stack[0][2] ),
    .I2(\stack[1][2] ),
    .I3(\stack[2][2] ),
    .S0(_00901_),
    .S1(_00902_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05358_ (.I(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05359_ (.I0(\stack[7][2] ),
    .I1(\stack[4][2] ),
    .I2(\stack[5][2] ),
    .I3(\stack[6][2] ),
    .S0(_00811_),
    .S1(_00891_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05360_ (.A1(_00894_),
    .A2(_00905_),
    .B(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05361_ (.A1(_00889_),
    .A2(_00911_),
    .B(_00913_),
    .C(_00878_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05362_ (.A1(_00781_),
    .A2(_00909_),
    .A3(_00914_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05363_ (.A1(_00898_),
    .A2(_00915_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05364_ (.I(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05365_ (.I(_00917_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05366_ (.I(_00918_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05367_ (.I(_00919_),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05368_ (.I(_00908_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05369_ (.I(_00887_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05370_ (.I(_00921_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05371_ (.A1(_00883_),
    .A2(_00832_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05372_ (.I(_00923_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05373_ (.I(_00924_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05374_ (.I(_00881_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05375_ (.I(_00926_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05376_ (.I(_00902_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05377_ (.A1(_00927_),
    .A2(\stack[0][3] ),
    .B1(\stack[1][3] ),
    .B2(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05378_ (.A1(_00925_),
    .A2(_00929_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05379_ (.I(_00786_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05380_ (.I(_00931_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05381_ (.I(_00923_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05382_ (.I(_00933_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05383_ (.A1(_00932_),
    .A2(\stack[3][3] ),
    .B1(_00934_),
    .B2(\stack[2][3] ),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05384_ (.A1(_00922_),
    .A2(_00930_),
    .A3(_00935_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05385_ (.I(_00799_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05386_ (.I(_00937_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05387_ (.A1(\stack[6][3] ),
    .A2(_00934_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05388_ (.I(_00790_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05389_ (.I(_00940_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05390_ (.I(_00941_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05391_ (.I0(\stack[5][3] ),
    .I1(\stack[4][3] ),
    .S(_00942_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05392_ (.I(_00883_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05393_ (.I(_00801_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05394_ (.A1(_00944_),
    .A2(_00945_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05395_ (.A1(\stack[7][3] ),
    .A2(_00905_),
    .B1(_00943_),
    .B2(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05396_ (.A1(_00938_),
    .A2(_00939_),
    .A3(_00947_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05397_ (.A1(_00920_),
    .A2(_00936_),
    .A3(_00948_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05398_ (.I(_00781_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05399_ (.I0(\stack[11][3] ),
    .I1(\stack[8][3] ),
    .I2(\stack[9][3] ),
    .I3(\stack[10][3] ),
    .S0(_00942_),
    .S1(_00928_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05400_ (.I(_00951_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05401_ (.I(_00926_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05402_ (.I(_00884_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05403_ (.I0(\stack[15][3] ),
    .I1(\stack[12][3] ),
    .I2(\stack[13][3] ),
    .I3(\stack[14][3] ),
    .S0(_00953_),
    .S1(_00954_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05404_ (.A1(_00894_),
    .A2(_00905_),
    .B(_00955_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05405_ (.A1(_00922_),
    .A2(_00952_),
    .B(_00956_),
    .C(_00908_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05406_ (.A1(_00950_),
    .A2(_00957_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05407_ (.I(_00772_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05408_ (.I(_00959_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05409_ (.I(_00887_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05410_ (.I(_00847_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05411_ (.I(_00962_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05412_ (.A1(_00927_),
    .A2(\stack[20][3] ),
    .B1(\stack[21][3] ),
    .B2(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05413_ (.A1(_00963_),
    .A2(_00927_),
    .A3(\stack[22][3] ),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05414_ (.A1(_00934_),
    .A2(_00964_),
    .B(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05415_ (.A1(\stack[23][3] ),
    .A2(_00960_),
    .B(_00961_),
    .C(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05416_ (.I(_00945_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05417_ (.I(_00962_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05418_ (.I0(\stack[19][3] ),
    .I1(\stack[16][3] ),
    .I2(\stack[17][3] ),
    .I3(\stack[18][3] ),
    .S0(_00968_),
    .S1(_00969_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05419_ (.A1(_00938_),
    .A2(_00970_),
    .B(_00908_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05420_ (.I(_00799_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05421_ (.I0(\stack[27][3] ),
    .I1(\stack[24][3] ),
    .I2(\stack[25][3] ),
    .I3(\stack[26][3] ),
    .S0(_00968_),
    .S1(_00963_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05422_ (.I(_00878_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05423_ (.A1(_00972_),
    .A2(_00973_),
    .B(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05424_ (.I0(\stack[31][3] ),
    .I1(\stack[28][3] ),
    .I2(\stack[29][3] ),
    .I3(\stack[30][3] ),
    .S0(_00968_),
    .S1(_00963_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05425_ (.A1(_00922_),
    .A2(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05426_ (.A1(_00967_),
    .A2(_00971_),
    .B1(_00975_),
    .B2(_00977_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05427_ (.I(_00854_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05428_ (.A1(_00949_),
    .A2(_00958_),
    .B1(_00978_),
    .B2(_00979_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05429_ (.I(_00980_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05430_ (.I(_00981_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05431_ (.I(_00982_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05432_ (.I(_00983_),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05433_ (.I(_00923_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05434_ (.A1(_00968_),
    .A2(\stack[4][4] ),
    .B1(\stack[5][4] ),
    .B2(_00928_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05435_ (.A1(_00984_),
    .A2(_00985_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05436_ (.A1(\stack[6][4] ),
    .A2(_00984_),
    .B1(_00959_),
    .B2(\stack[7][4] ),
    .C(_00921_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05437_ (.A1(_00945_),
    .A2(\stack[0][4] ),
    .B1(\stack[1][4] ),
    .B2(_00944_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05438_ (.A1(_00923_),
    .A2(_00988_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05439_ (.A1(_00931_),
    .A2(\stack[3][4] ),
    .B1(_00924_),
    .B2(\stack[2][4] ),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05440_ (.A1(_00889_),
    .A2(_00989_),
    .A3(_00990_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05441_ (.A1(_00986_),
    .A2(_00987_),
    .B(_00991_),
    .C(_00879_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05442_ (.I(_00959_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05443_ (.A1(\stack[15][4] ),
    .A2(_00993_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05444_ (.I0(\stack[13][4] ),
    .I1(\stack[12][4] ),
    .S(_00942_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05445_ (.A1(\stack[14][4] ),
    .A2(_00925_),
    .B1(_00946_),
    .B2(_00995_),
    .C(_00921_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05446_ (.I0(\stack[11][4] ),
    .I1(\stack[8][4] ),
    .I2(\stack[9][4] ),
    .I3(\stack[10][4] ),
    .S0(_00953_),
    .S1(_00954_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05447_ (.A1(_00937_),
    .A2(_00997_),
    .B(_00879_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05448_ (.A1(_00994_),
    .A2(_00996_),
    .B(_00998_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05449_ (.A1(_00950_),
    .A2(_00992_),
    .A3(_00999_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05450_ (.A1(_00942_),
    .A2(\stack[20][4] ),
    .B1(\stack[21][4] ),
    .B2(_00962_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05451_ (.A1(_00933_),
    .A2(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05452_ (.A1(\stack[22][4] ),
    .A2(_00984_),
    .B1(_00993_),
    .B2(\stack[23][4] ),
    .C(_01002_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05453_ (.A1(_00945_),
    .A2(\stack[16][4] ),
    .B1(\stack[17][4] ),
    .B2(_00962_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05454_ (.A1(_00924_),
    .A2(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05455_ (.A1(_00931_),
    .A2(\stack[19][4] ),
    .B1(_00933_),
    .B2(\stack[18][4] ),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05456_ (.A1(_00921_),
    .A2(_01005_),
    .A3(_01006_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05457_ (.A1(_00972_),
    .A2(_01003_),
    .B(_01007_),
    .C(_00974_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05458_ (.A1(_00924_),
    .A2(_00959_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05459_ (.I(_00767_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05460_ (.I(_01010_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05461_ (.I(_01011_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05462_ (.I(_00855_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05463_ (.I(_01013_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05464_ (.I(_01014_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05465_ (.A1(_01012_),
    .A2(\stack[28][4] ),
    .B1(\stack[29][4] ),
    .B2(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05466_ (.A1(_01009_),
    .A2(_01016_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05467_ (.A1(\stack[30][4] ),
    .A2(_00925_),
    .B1(_00993_),
    .B2(\stack[31][4] ),
    .C(_00961_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05468_ (.I0(\stack[27][4] ),
    .I1(\stack[24][4] ),
    .I2(\stack[25][4] ),
    .I3(\stack[26][4] ),
    .S0(_00953_),
    .S1(_00954_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05469_ (.A1(_00937_),
    .A2(_01019_),
    .B(_00879_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05470_ (.A1(_01017_),
    .A2(_01018_),
    .B(_01020_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05471_ (.A1(_00854_),
    .A2(_01008_),
    .A3(_01021_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05472_ (.A1(_01000_),
    .A2(_01022_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05473_ (.I(_01023_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05474_ (.I(_01024_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05475_ (.I(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05476_ (.I(_01026_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05477_ (.I(_01027_),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05478_ (.I(_00961_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05479_ (.I(_00953_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05480_ (.I(_01029_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05481_ (.I(_00928_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05482_ (.I0(\stack[23][5] ),
    .I1(\stack[20][5] ),
    .I2(\stack[21][5] ),
    .I3(\stack[22][5] ),
    .S0(_01030_),
    .S1(_01031_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05483_ (.I(_00925_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05484_ (.A1(_01030_),
    .A2(\stack[16][5] ),
    .B1(\stack[17][5] ),
    .B2(_01031_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05485_ (.A1(_01033_),
    .A2(_01034_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05486_ (.I(_00932_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05487_ (.A1(_01036_),
    .A2(\stack[19][5] ),
    .B1(_01033_),
    .B2(\stack[18][5] ),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05488_ (.A1(_01028_),
    .A2(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05489_ (.A1(_01028_),
    .A2(_01032_),
    .B1(_01035_),
    .B2(_01038_),
    .C(_00920_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05490_ (.I(_00972_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05491_ (.I(_01009_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05492_ (.I(_01012_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05493_ (.I(_01015_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05494_ (.A1(_01042_),
    .A2(\stack[24][5] ),
    .B1(\stack[25][5] ),
    .B2(_01043_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05495_ (.I(_00984_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05496_ (.A1(\stack[26][5] ),
    .A2(_01045_),
    .B1(_00960_),
    .B2(\stack[27][5] ),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05497_ (.A1(_01041_),
    .A2(_01044_),
    .B(_01046_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05498_ (.A1(_01042_),
    .A2(\stack[28][5] ),
    .B1(\stack[29][5] ),
    .B2(_01043_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05499_ (.I(_00933_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05500_ (.A1(\stack[30][5] ),
    .A2(_01049_),
    .B1(_00960_),
    .B2(\stack[31][5] ),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05501_ (.I(_00937_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05502_ (.A1(_01009_),
    .A2(_01048_),
    .B(_01050_),
    .C(_01051_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05503_ (.I(_00974_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05504_ (.A1(_01040_),
    .A2(_01047_),
    .B(_01052_),
    .C(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05505_ (.A1(_01039_),
    .A2(_01054_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05506_ (.A1(_01030_),
    .A2(\stack[0][5] ),
    .B1(\stack[1][5] ),
    .B2(_01031_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05507_ (.A1(_01049_),
    .A2(_01056_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05508_ (.A1(_01036_),
    .A2(\stack[3][5] ),
    .B1(_01045_),
    .B2(\stack[2][5] ),
    .C(_00972_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05509_ (.I0(\stack[7][5] ),
    .I1(\stack[4][5] ),
    .I2(\stack[5][5] ),
    .I3(\stack[6][5] ),
    .S0(_01029_),
    .S1(_00969_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05510_ (.A1(_00922_),
    .A2(_01059_),
    .B(_00920_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05511_ (.A1(_01057_),
    .A2(_01058_),
    .B(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05512_ (.I(_00993_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05513_ (.A1(\stack[15][5] ),
    .A2(_01062_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05514_ (.I(_00946_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05515_ (.I0(\stack[13][5] ),
    .I1(\stack[12][5] ),
    .S(_00927_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05516_ (.A1(\stack[14][5] ),
    .A2(_01045_),
    .B1(_01064_),
    .B2(_01065_),
    .C(_00961_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05517_ (.I0(\stack[11][5] ),
    .I1(\stack[8][5] ),
    .I2(\stack[9][5] ),
    .I3(\stack[10][5] ),
    .S0(_01029_),
    .S1(_00969_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05518_ (.A1(_00938_),
    .A2(_01067_),
    .B(_00974_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05519_ (.A1(_01063_),
    .A2(_01066_),
    .B(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05520_ (.A1(_01061_),
    .A2(_01069_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05521_ (.A1(_00979_),
    .A2(_01070_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05522_ (.A1(_00979_),
    .A2(_01055_),
    .B(_01071_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05523_ (.I(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05524_ (.I(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05525_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05526_ (.I(_01075_),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05527_ (.I(_00960_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05528_ (.I(_01042_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05529_ (.I(_01043_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05530_ (.A1(_01077_),
    .A2(\stack[12][6] ),
    .B1(\stack[13][6] ),
    .B2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05531_ (.I(_01049_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05532_ (.A1(\stack[14][6] ),
    .A2(_01080_),
    .B1(_01076_),
    .B2(\stack[15][6] ),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05533_ (.A1(_01076_),
    .A2(_01079_),
    .B(_01081_),
    .C(_01040_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05534_ (.I(_01012_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05535_ (.I(_01015_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05536_ (.A1(_01083_),
    .A2(\stack[8][6] ),
    .B1(\stack[9][6] ),
    .B2(_01084_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05537_ (.A1(_01062_),
    .A2(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05538_ (.I(_00932_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05539_ (.A1(_01087_),
    .A2(\stack[11][6] ),
    .B1(_01080_),
    .B2(\stack[10][6] ),
    .C(_01040_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05540_ (.I(_00920_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05541_ (.A1(_01086_),
    .A2(_01088_),
    .B(_01089_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05542_ (.A1(_01042_),
    .A2(\stack[0][6] ),
    .B1(\stack[1][6] ),
    .B2(_01084_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05543_ (.A1(_01041_),
    .A2(_01091_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05544_ (.I(_00932_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05545_ (.I(_00934_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05546_ (.A1(_01093_),
    .A2(\stack[3][6] ),
    .B1(_01094_),
    .B2(\stack[2][6] ),
    .C(_01051_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05547_ (.A1(_01012_),
    .A2(\stack[4][6] ),
    .B1(\stack[5][6] ),
    .B2(_01043_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05548_ (.A1(\stack[6][6] ),
    .A2(_01049_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05549_ (.A1(_01009_),
    .A2(_01096_),
    .B(_01097_),
    .C(_00938_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05550_ (.A1(\stack[7][6] ),
    .A2(_01062_),
    .B(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05551_ (.A1(_01092_),
    .A2(_01095_),
    .B(_01099_),
    .C(_01053_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05552_ (.A1(_01082_),
    .A2(_01090_),
    .B(_01100_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05553_ (.I(_01028_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05554_ (.I(_01041_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05555_ (.A1(_01077_),
    .A2(\stack[28][6] ),
    .B1(\stack[29][6] ),
    .B2(_01078_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05556_ (.I(_01045_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05557_ (.A1(\stack[30][6] ),
    .A2(_01105_),
    .B1(_01076_),
    .B2(\stack[31][6] ),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05558_ (.A1(_01103_),
    .A2(_01104_),
    .B(_01106_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05559_ (.A1(_01083_),
    .A2(\stack[24][6] ),
    .B1(\stack[25][6] ),
    .B2(_01078_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05560_ (.A1(_01093_),
    .A2(\stack[27][6] ),
    .B1(_01094_),
    .B2(\stack[26][6] ),
    .C(_01051_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05561_ (.A1(_01103_),
    .A2(_01108_),
    .B(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05562_ (.A1(_01102_),
    .A2(_01107_),
    .B(_01110_),
    .C(_01053_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05563_ (.I0(\stack[23][6] ),
    .I1(\stack[20][6] ),
    .I2(\stack[21][6] ),
    .I3(\stack[22][6] ),
    .S0(_01030_),
    .S1(_01031_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05564_ (.I(_01029_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05565_ (.I(_00969_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05566_ (.A1(_01113_),
    .A2(\stack[16][6] ),
    .B1(\stack[17][6] ),
    .B2(_01114_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05567_ (.A1(_01094_),
    .A2(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05568_ (.A1(_01036_),
    .A2(\stack[19][6] ),
    .B1(_01033_),
    .B2(\stack[18][6] ),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05569_ (.A1(_01028_),
    .A2(_01117_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05570_ (.A1(_01102_),
    .A2(_01112_),
    .B1(_01116_),
    .B2(_01118_),
    .C(_01089_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05571_ (.A1(_00950_),
    .A2(_01119_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05572_ (.A1(_00979_),
    .A2(_01101_),
    .B1(_01111_),
    .B2(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05573_ (.I(_01121_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05574_ (.I(_01122_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05575_ (.I(_01123_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05576_ (.I(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05577_ (.I(_01125_),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05578_ (.I(_00950_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05579_ (.I(_01102_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05580_ (.I0(\stack[7][7] ),
    .I1(\stack[4][7] ),
    .I2(\stack[5][7] ),
    .I3(\stack[6][7] ),
    .S0(_01113_),
    .S1(_01114_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05581_ (.I(_01041_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05582_ (.I(_01083_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05583_ (.I(_01084_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05584_ (.A1(_01130_),
    .A2(\stack[0][7] ),
    .B1(\stack[1][7] ),
    .B2(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05585_ (.I(_01093_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05586_ (.I(_01051_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05587_ (.A1(_01133_),
    .A2(\stack[3][7] ),
    .B1(_01105_),
    .B2(\stack[2][7] ),
    .C(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05588_ (.A1(_01129_),
    .A2(_01132_),
    .B(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05589_ (.I(_01089_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05590_ (.A1(_01127_),
    .A2(_01128_),
    .B(_01136_),
    .C(_01137_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05591_ (.A1(_01130_),
    .A2(\stack[12][7] ),
    .B1(\stack[13][7] ),
    .B2(_01131_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05592_ (.I(_01094_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05593_ (.I(_01062_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05594_ (.A1(\stack[14][7] ),
    .A2(_01140_),
    .B1(_01141_),
    .B2(\stack[15][7] ),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05595_ (.A1(_01129_),
    .A2(_01139_),
    .B(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05596_ (.I(_01083_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05597_ (.A1(_01144_),
    .A2(\stack[8][7] ),
    .B1(\stack[9][7] ),
    .B2(_01131_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05598_ (.A1(_01087_),
    .A2(\stack[11][7] ),
    .B1(_01105_),
    .B2(\stack[10][7] ),
    .C(_01040_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05599_ (.A1(_01129_),
    .A2(_01145_),
    .B(_01146_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05600_ (.A1(_01127_),
    .A2(_01143_),
    .B(_01147_),
    .C(_01053_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05601_ (.A1(_01138_),
    .A2(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05602_ (.I(_01084_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05603_ (.A1(_01144_),
    .A2(\stack[16][7] ),
    .B1(\stack[17][7] ),
    .B2(_01150_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05604_ (.A1(\stack[18][7] ),
    .A2(_01140_),
    .B1(_01141_),
    .B2(\stack[19][7] ),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05605_ (.A1(_01129_),
    .A2(_01151_),
    .B(_01152_),
    .C(_01127_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05606_ (.A1(_01077_),
    .A2(\stack[20][7] ),
    .B1(\stack[21][7] ),
    .B2(_01078_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05607_ (.A1(\stack[22][7] ),
    .A2(_01080_),
    .B1(_01076_),
    .B2(\stack[23][7] ),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05608_ (.A1(_01103_),
    .A2(_01154_),
    .B(_01155_),
    .C(_01134_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05609_ (.A1(_01137_),
    .A2(_01156_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05610_ (.A1(_01144_),
    .A2(\stack[28][7] ),
    .B1(\stack[29][7] ),
    .B2(_01150_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05611_ (.A1(\stack[30][7] ),
    .A2(_01140_),
    .B1(_01141_),
    .B2(\stack[31][7] ),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05612_ (.A1(_01141_),
    .A2(_01158_),
    .B(_01159_),
    .C(_01134_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05613_ (.A1(_01077_),
    .A2(\stack[24][7] ),
    .B1(\stack[25][7] ),
    .B2(_01150_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05614_ (.A1(_01103_),
    .A2(_01161_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05615_ (.A1(_01133_),
    .A2(\stack[27][7] ),
    .B1(_01140_),
    .B2(\stack[26][7] ),
    .C(_01134_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05616_ (.A1(_01162_),
    .A2(_01163_),
    .B(_01137_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05617_ (.A1(_01153_),
    .A2(_01157_),
    .B1(_01160_),
    .B2(_01164_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05618_ (.A1(_01126_),
    .A2(_01165_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05619_ (.A1(_01126_),
    .A2(_01149_),
    .B(_01166_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05620_ (.I(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05621_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05622_ (.I(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05623_ (.I(_01170_),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05624_ (.I(\mem.select ),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05625_ (.I(\mem.sram_enable ),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05626_ (.I(net188),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05627_ (.A1(net190),
    .A2(net189),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05628_ (.A1(_01173_),
    .A2(_01174_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05629_ (.A1(\mem.mem_dff.memory_type_data ),
    .A2(_01175_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05630_ (.A1(net189),
    .A2(net188),
    .B(_01176_),
    .C(net190),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05631_ (.A1(_01171_),
    .A2(_01172_),
    .A3(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05632_ (.I(_01178_),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05633_ (.A1(\intr_enable[0] ),
    .A2(\intr[0] ),
    .B1(\intr[1] ),
    .B2(\intr_enable[1] ),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05634_ (.A1(edge_interrupts),
    .A2(prev_level_interrupt),
    .B(_01179_),
    .ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05635_ (.A1(wb_write_ack),
    .A2(wb_read_ack),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05636_ (.I(_01180_),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05637_ (.I(_00839_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05638_ (.I(_01181_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05639_ (.I(_01182_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05640_ (.I(net132),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05641_ (.I(net131),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05642_ (.I(_01185_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05643_ (.A1(net134),
    .A2(net133),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05644_ (.A1(_01184_),
    .A2(_01186_),
    .A3(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05645_ (.I(_01188_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05646_ (.I(net130),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05647_ (.I(_01190_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05648_ (.I(net129),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05649_ (.A1(net258),
    .A2(net158),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05650_ (.A1(_01191_),
    .A2(_01192_),
    .A3(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05651_ (.A1(_01189_),
    .A2(_01194_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05652_ (.I(net258),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05653_ (.I(net158),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05654_ (.A1(_01196_),
    .A2(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05655_ (.A1(_01190_),
    .A2(_01192_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05656_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05657_ (.A1(_01184_),
    .A2(_01185_),
    .A3(_01187_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05658_ (.I(_01201_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05659_ (.A1(_01198_),
    .A2(_01200_),
    .A3(_01202_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05660_ (.A1(_01195_),
    .A2(_01203_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05661_ (.A1(_01188_),
    .A2(_01198_),
    .A3(_01200_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05662_ (.A1(net258),
    .A2(_01197_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05663_ (.I(_01192_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05664_ (.A1(_01190_),
    .A2(_01207_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05665_ (.A1(_01189_),
    .A2(_01206_),
    .A3(_01208_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05666_ (.A1(_01205_),
    .A2(_01209_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05667_ (.I(net159),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05668_ (.I(net158),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05669_ (.A1(_01211_),
    .A2(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05670_ (.I(_01184_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05671_ (.I(_01185_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05672_ (.I(net134),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05673_ (.I(net133),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05674_ (.I(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05675_ (.A1(_01216_),
    .A2(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05676_ (.A1(_01214_),
    .A2(_01215_),
    .A3(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05677_ (.A1(_01200_),
    .A2(_01213_),
    .A3(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05678_ (.I(net134),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05679_ (.A1(_01222_),
    .A2(net133),
    .A3(net132),
    .A4(net131),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05680_ (.I(_01223_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05681_ (.A1(_01224_),
    .A2(_01194_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05682_ (.A1(_01221_),
    .A2(_01225_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05683_ (.I(_01190_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05684_ (.I(_01192_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05685_ (.A1(_01227_),
    .A2(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05686_ (.A1(_01189_),
    .A2(_01229_),
    .A3(_01213_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05687_ (.A1(_01204_),
    .A2(_01210_),
    .A3(_01226_),
    .A4(_01230_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05688_ (.I(_01231_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05689_ (.I(_01184_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05690_ (.A1(_01233_),
    .A2(_01215_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05691_ (.A1(net130),
    .A2(net129),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05692_ (.A1(_01193_),
    .A2(_01234_),
    .A3(_01219_),
    .A4(_01235_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05693_ (.A1(_01188_),
    .A2(_01198_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05694_ (.A1(_01224_),
    .A2(_01206_),
    .A3(_01229_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05695_ (.A1(_01235_),
    .A2(_01237_),
    .B(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05696_ (.I(_01239_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05697_ (.A1(_01223_),
    .A2(_01213_),
    .A3(_01208_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05698_ (.A1(_01216_),
    .A2(_01217_),
    .A3(_01233_),
    .A4(_01185_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05699_ (.A1(_01206_),
    .A2(_01199_),
    .A3(_01242_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05700_ (.A1(_01241_),
    .A2(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05701_ (.A1(_01211_),
    .A2(_01212_),
    .A3(_01235_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _05702_ (.A1(_01206_),
    .A2(_01199_),
    .A3(_01201_),
    .B1(_01245_),
    .B2(_01223_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05703_ (.A1(_01199_),
    .A2(_01201_),
    .A3(_01213_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05704_ (.A1(_01194_),
    .A2(_01201_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05705_ (.A1(_01246_),
    .A2(_01247_),
    .A3(_01248_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05706_ (.A1(_01224_),
    .A2(_01208_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05707_ (.A1(_01193_),
    .A2(_01250_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05708_ (.A1(_01244_),
    .A2(_01249_),
    .A3(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05709_ (.A1(_01236_),
    .A2(_01240_),
    .A3(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05710_ (.A1(_01232_),
    .A2(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05711_ (.I(_00773_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05712_ (.A1(_01255_),
    .A2(_01087_),
    .A3(_01105_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05713_ (.A1(_00778_),
    .A2(_01256_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05714_ (.A1(_00774_),
    .A2(_00766_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05715_ (.I(_01258_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05716_ (.I(_01259_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05717_ (.I(_00881_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05718_ (.I0(\stack[2][2] ),
    .I1(\stack[3][2] ),
    .I2(\stack[0][2] ),
    .I3(\stack[1][2] ),
    .S0(_01261_),
    .S1(_00902_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05719_ (.A1(_00941_),
    .A2(\stack[5][2] ),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05720_ (.I(_01014_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05721_ (.A1(_00774_),
    .A2(_00766_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05722_ (.I(_01265_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05723_ (.I(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05724_ (.A1(_01264_),
    .A2(\stack[4][2] ),
    .B(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05725_ (.A1(_01264_),
    .A2(\stack[6][2] ),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05726_ (.A1(net137),
    .A2(_00775_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05727_ (.I(_01270_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05728_ (.I(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05729_ (.A1(_00941_),
    .A2(\stack[7][2] ),
    .B(_01272_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05730_ (.A1(_00805_),
    .A2(_01270_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05731_ (.I(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05732_ (.A1(_01263_),
    .A2(_01268_),
    .B1(_01269_),
    .B2(_01273_),
    .C(_01275_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05733_ (.A1(_01260_),
    .A2(_01262_),
    .B(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05734_ (.I(_01274_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05735_ (.I(_01278_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05736_ (.I(_01270_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05737_ (.A1(_01280_),
    .A2(_01265_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05738_ (.I(_01281_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05739_ (.I0(\stack[10][2] ),
    .I1(\stack[11][2] ),
    .S(_00940_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05740_ (.I0(\stack[8][2] ),
    .I1(\stack[9][2] ),
    .S(_00857_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05741_ (.I(_00786_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05742_ (.I(_01285_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05743_ (.A1(_01011_),
    .A2(_01283_),
    .B1(_01284_),
    .B2(_01286_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05744_ (.I0(\stack[12][2] ),
    .I1(\stack[13][2] ),
    .S(_00857_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05745_ (.I0(\stack[14][2] ),
    .I1(\stack[15][2] ),
    .S(_00900_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05746_ (.I(_01280_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05747_ (.I(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05748_ (.A1(_01267_),
    .A2(_01288_),
    .B1(_01289_),
    .B2(_01291_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05749_ (.A1(_01282_),
    .A2(_01287_),
    .B(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05750_ (.A1(_01279_),
    .A2(_01293_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(_01277_),
    .A2(_01294_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05752_ (.I0(\stack[18][2] ),
    .I1(\stack[19][2] ),
    .I2(\stack[16][2] ),
    .I3(\stack[17][2] ),
    .S0(_00792_),
    .S1(_00884_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05753_ (.A1(_01260_),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05754_ (.I(_01280_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05755_ (.I(_01298_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05756_ (.I0(\stack[22][2] ),
    .I1(\stack[23][2] ),
    .S(_01261_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05757_ (.I0(\stack[20][2] ),
    .I1(\stack[21][2] ),
    .S(_00901_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05758_ (.I(_01265_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05759_ (.I(_01302_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05760_ (.I(_01303_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05761_ (.A1(_00773_),
    .A2(_01270_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05762_ (.I(_01305_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05763_ (.I(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05764_ (.A1(_01299_),
    .A2(_01300_),
    .B1(_01301_),
    .B2(_01304_),
    .C(_01307_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05765_ (.I0(\stack[24][2] ),
    .I1(\stack[25][2] ),
    .S(_00901_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05766_ (.A1(_01264_),
    .A2(\stack[26][2] ),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05767_ (.A1(_00926_),
    .A2(\stack[27][2] ),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05768_ (.A1(_01310_),
    .A2(_01311_),
    .B(_00944_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05769_ (.I(_01258_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05770_ (.A1(_00954_),
    .A2(_01309_),
    .B(_01312_),
    .C(_01313_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05771_ (.I(\stack[31][2] ),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05772_ (.A1(_01264_),
    .A2(\stack[30][2] ),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05773_ (.A1(_01015_),
    .A2(_01315_),
    .B(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05774_ (.I0(\stack[28][2] ),
    .I1(\stack[29][2] ),
    .S(_00882_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05775_ (.A1(_01299_),
    .A2(_01317_),
    .B1(_01318_),
    .B2(_01304_),
    .C(_01279_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05776_ (.A1(_01297_),
    .A2(_01308_),
    .B1(_01314_),
    .B2(_01319_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05777_ (.I(_00851_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05778_ (.I0(_01295_),
    .I1(_01320_),
    .S(_01321_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05779_ (.I0(\stack[26][0] ),
    .I1(\stack[27][0] ),
    .S(_00792_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05780_ (.I0(\stack[24][0] ),
    .I1(\stack[25][0] ),
    .S(_00792_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05781_ (.A1(_01011_),
    .A2(_01323_),
    .B1(_01324_),
    .B2(_01286_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05782_ (.I(\stack[31][0] ),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05783_ (.A1(_01261_),
    .A2(\stack[30][0] ),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05784_ (.A1(_00941_),
    .A2(_01326_),
    .B(_01327_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05785_ (.I(_00899_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05786_ (.I(_01329_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05787_ (.I0(\stack[28][0] ),
    .I1(\stack[29][0] ),
    .S(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05788_ (.A1(_01299_),
    .A2(_01328_),
    .B1(_01331_),
    .B2(_01304_),
    .C(_01275_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05789_ (.A1(_01282_),
    .A2(_01325_),
    .B(_01332_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05790_ (.I0(\stack[18][0] ),
    .I1(\stack[19][0] ),
    .I2(\stack[16][0] ),
    .I3(\stack[17][0] ),
    .S0(_01330_),
    .S1(_00844_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05791_ (.A1(_01260_),
    .A2(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05792_ (.I0(\stack[22][0] ),
    .I1(\stack[23][0] ),
    .S(_00882_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05793_ (.I0(\stack[20][0] ),
    .I1(\stack[21][0] ),
    .S(_00811_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05794_ (.A1(_01299_),
    .A2(_01336_),
    .B1(_01337_),
    .B2(_01304_),
    .C(_01307_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05795_ (.A1(_01335_),
    .A2(_01338_),
    .B(_01321_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05796_ (.I0(\stack[4][0] ),
    .I1(\stack[5][0] ),
    .S(_00843_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05797_ (.I0(\stack[6][0] ),
    .I1(\stack[7][0] ),
    .S(_00801_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05798_ (.I(_01290_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05799_ (.I0(\stack[2][0] ),
    .I1(\stack[3][0] ),
    .I2(\stack[0][0] ),
    .I3(\stack[1][0] ),
    .S0(_00790_),
    .S1(_00802_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05800_ (.A1(_01258_),
    .A2(_01343_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05801_ (.A1(_01267_),
    .A2(_01340_),
    .B1(_01341_),
    .B2(_01342_),
    .C(_01344_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05802_ (.I0(\stack[8][0] ),
    .I1(\stack[9][0] ),
    .S(_00822_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05803_ (.I(\stack[11][0] ),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05804_ (.A1(_00832_),
    .A2(\stack[10][0] ),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05805_ (.A1(_01261_),
    .A2(_01347_),
    .B(_01348_),
    .C(_00844_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05806_ (.A1(_00944_),
    .A2(_01346_),
    .B(_01349_),
    .C(_01313_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05807_ (.I0(\stack[12][0] ),
    .I1(\stack[13][0] ),
    .S(_01330_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05808_ (.I(\stack[15][0] ),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05809_ (.A1(_01330_),
    .A2(\stack[14][0] ),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05810_ (.A1(_00926_),
    .A2(_01352_),
    .B(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05811_ (.I(_01274_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05812_ (.A1(_01267_),
    .A2(_01351_),
    .B1(_01354_),
    .B2(_01342_),
    .C(_01355_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05813_ (.I(_00777_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05814_ (.A1(_01279_),
    .A2(_01345_),
    .B1(_01350_),
    .B2(_01356_),
    .C(_01357_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05815_ (.A1(_01333_),
    .A2(_01339_),
    .B(_01358_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05816_ (.I(_00769_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05817_ (.I0(\stack[18][7] ),
    .I1(\stack[19][7] ),
    .S(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05818_ (.I0(\stack[16][7] ),
    .I1(\stack[17][7] ),
    .S(_01013_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05819_ (.I(_00786_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05820_ (.A1(_00803_),
    .A2(_01361_),
    .B1(_01362_),
    .B2(_01363_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05821_ (.I0(\stack[20][7] ),
    .I1(\stack[21][7] ),
    .S(_01360_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05822_ (.I0(\stack[22][7] ),
    .I1(\stack[23][7] ),
    .S(_01013_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05823_ (.A1(_01303_),
    .A2(_01365_),
    .B1(_01366_),
    .B2(_01290_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05824_ (.A1(_01291_),
    .A2(_01364_),
    .B(_01278_),
    .C(_01367_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05825_ (.I(_00820_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05826_ (.I0(\stack[24][7] ),
    .I1(\stack[25][7] ),
    .S(_01369_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05827_ (.I(_00855_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05828_ (.I0(\stack[26][7] ),
    .I1(\stack[27][7] ),
    .S(_01371_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05829_ (.A1(_01363_),
    .A2(_01370_),
    .B1(_01372_),
    .B2(_00803_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05830_ (.I(_00820_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05831_ (.I0(\stack[28][7] ),
    .I1(\stack[29][7] ),
    .S(_01374_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05832_ (.I0(\stack[30][7] ),
    .I1(\stack[31][7] ),
    .S(_01371_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05833_ (.A1(_01303_),
    .A2(_01375_),
    .B1(_01376_),
    .B2(_01298_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05834_ (.A1(_01291_),
    .A2(_01373_),
    .B(_01377_),
    .C(_01306_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05835_ (.A1(_01368_),
    .A2(_01378_),
    .B(_00852_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05836_ (.I(_01281_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05837_ (.I0(\stack[10][7] ),
    .I1(\stack[11][7] ),
    .S(_00868_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05838_ (.I0(\stack[8][7] ),
    .I1(\stack[9][7] ),
    .S(_00800_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05839_ (.A1(_01010_),
    .A2(_01381_),
    .B1(_01382_),
    .B2(_01285_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05840_ (.I0(\stack[12][7] ),
    .I1(\stack[13][7] ),
    .S(_00770_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05841_ (.I0(\stack[14][7] ),
    .I1(\stack[15][7] ),
    .S(_01013_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05842_ (.A1(_01266_),
    .A2(_01384_),
    .B1(_01385_),
    .B2(_01290_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05843_ (.A1(_01380_),
    .A2(_01383_),
    .B(_01386_),
    .C(_01306_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05844_ (.I0(\stack[2][7] ),
    .I1(\stack[3][7] ),
    .I2(\stack[0][7] ),
    .I3(\stack[1][7] ),
    .S0(_00856_),
    .S1(_00869_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05845_ (.A1(_01259_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05846_ (.I(_01266_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05847_ (.I(_00899_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05848_ (.I0(\stack[4][7] ),
    .I1(\stack[5][7] ),
    .S(_01391_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05849_ (.I0(\stack[6][7] ),
    .I1(\stack[7][7] ),
    .S(_01369_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05850_ (.I(_01271_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05851_ (.A1(_01390_),
    .A2(_01392_),
    .B1(_01393_),
    .B2(_01394_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05852_ (.A1(_01278_),
    .A2(_01389_),
    .A3(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05853_ (.A1(_01387_),
    .A2(_01396_),
    .B(_00777_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05854_ (.I(_01258_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05855_ (.I0(\stack[18][6] ),
    .I1(\stack[19][6] ),
    .I2(\stack[16][6] ),
    .I3(\stack[17][6] ),
    .S0(_00868_),
    .S1(_00890_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05856_ (.A1(_01398_),
    .A2(_01399_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05857_ (.I(_01266_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05858_ (.I0(\stack[20][6] ),
    .I1(\stack[21][6] ),
    .S(_00810_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05859_ (.I(_00809_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05860_ (.I0(\stack[22][6] ),
    .I1(\stack[23][6] ),
    .S(_01403_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05861_ (.I(_01271_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05862_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01404_),
    .B2(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05863_ (.A1(_01355_),
    .A2(_01400_),
    .A3(_01406_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05864_ (.I(_01281_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05865_ (.I(_01010_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05866_ (.I(_00880_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05867_ (.I0(\stack[26][6] ),
    .I1(\stack[27][6] ),
    .S(_01410_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05868_ (.I(_00809_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05869_ (.I0(\stack[24][6] ),
    .I1(\stack[25][6] ),
    .S(_01412_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05870_ (.I(_01285_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05871_ (.A1(_01409_),
    .A2(_01411_),
    .B1(_01413_),
    .B2(_01414_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05872_ (.I(_01302_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05873_ (.I(_00809_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05874_ (.I0(\stack[28][6] ),
    .I1(\stack[29][6] ),
    .S(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05875_ (.I0(\stack[30][6] ),
    .I1(\stack[31][6] ),
    .S(_01360_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05876_ (.I(_01271_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05877_ (.A1(_01416_),
    .A2(_01418_),
    .B1(_01419_),
    .B2(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05878_ (.I(_01306_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05879_ (.A1(_01408_),
    .A2(_01415_),
    .B(_01421_),
    .C(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05880_ (.I(_00852_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05881_ (.A1(_01407_),
    .A2(_01423_),
    .B(_01424_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05882_ (.I(_01010_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05883_ (.I(_00880_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05884_ (.I0(\stack[10][6] ),
    .I1(\stack[11][6] ),
    .S(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05885_ (.I0(\stack[8][6] ),
    .I1(\stack[9][6] ),
    .S(_01403_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05886_ (.I(_01285_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05887_ (.A1(_01426_),
    .A2(_01428_),
    .B1(_01429_),
    .B2(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05888_ (.I0(\stack[12][6] ),
    .I1(\stack[13][6] ),
    .S(_01412_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05889_ (.I0(\stack[14][6] ),
    .I1(\stack[15][6] ),
    .S(_00827_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05890_ (.I(_01280_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05891_ (.A1(_01416_),
    .A2(_01432_),
    .B1(_01433_),
    .B2(_01434_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05892_ (.I(_01305_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05893_ (.A1(_01408_),
    .A2(_01431_),
    .B(_01435_),
    .C(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05894_ (.I(_00820_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05895_ (.I0(\stack[2][6] ),
    .I1(\stack[3][6] ),
    .I2(\stack[0][6] ),
    .I3(\stack[1][6] ),
    .S0(_01438_),
    .S1(_00828_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05896_ (.A1(_01313_),
    .A2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05897_ (.I0(\stack[4][6] ),
    .I1(\stack[5][6] ),
    .S(_00881_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05898_ (.I(_00790_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05899_ (.I0(\stack[6][6] ),
    .I1(\stack[7][6] ),
    .S(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05900_ (.A1(_01401_),
    .A2(_01441_),
    .B1(_01443_),
    .B2(_01272_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05901_ (.A1(_01275_),
    .A2(_01440_),
    .A3(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05902_ (.I(_00777_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05903_ (.A1(_01437_),
    .A2(_01445_),
    .B(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05904_ (.A1(_01379_),
    .A2(_01397_),
    .A3(_01425_),
    .A4(_01447_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05905_ (.I0(\stack[18][3] ),
    .I1(\stack[19][3] ),
    .I2(\stack[16][3] ),
    .I3(\stack[17][3] ),
    .S0(_00800_),
    .S1(_00890_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05906_ (.A1(_01398_),
    .A2(_01449_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05907_ (.I0(\stack[20][3] ),
    .I1(\stack[21][3] ),
    .S(_00791_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05908_ (.I0(\stack[22][3] ),
    .I1(\stack[23][3] ),
    .S(_01403_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05909_ (.A1(_01401_),
    .A2(_01451_),
    .B1(_01452_),
    .B2(_01405_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05910_ (.A1(_01355_),
    .A2(_01450_),
    .A3(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05911_ (.I0(\stack[26][3] ),
    .I1(\stack[27][3] ),
    .S(_01410_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05912_ (.I0(\stack[24][3] ),
    .I1(\stack[25][3] ),
    .S(_01412_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05913_ (.A1(_01409_),
    .A2(_01455_),
    .B1(_01456_),
    .B2(_01414_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05914_ (.I0(\stack[28][3] ),
    .I1(\stack[29][3] ),
    .S(_01417_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05915_ (.I0(\stack[30][3] ),
    .I1(\stack[31][3] ),
    .S(_00821_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05916_ (.A1(_01416_),
    .A2(_01458_),
    .B1(_01459_),
    .B2(_01420_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05917_ (.A1(_01408_),
    .A2(_01457_),
    .B(_01460_),
    .C(_01422_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05918_ (.A1(_01454_),
    .A2(_01461_),
    .B(_01424_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05919_ (.I(_00880_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05920_ (.I0(\stack[10][3] ),
    .I1(\stack[11][3] ),
    .S(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05921_ (.I0(\stack[8][3] ),
    .I1(\stack[9][3] ),
    .S(_01427_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05922_ (.A1(_01426_),
    .A2(_01464_),
    .B1(_01465_),
    .B2(_01430_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05923_ (.I(_01302_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05924_ (.I0(\stack[12][3] ),
    .I1(\stack[13][3] ),
    .S(_01410_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05925_ (.I0(\stack[14][3] ),
    .I1(\stack[15][3] ),
    .S(_00770_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05926_ (.A1(_01467_),
    .A2(_01468_),
    .B1(_01469_),
    .B2(_01434_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05927_ (.A1(_01380_),
    .A2(_01466_),
    .B(_01470_),
    .C(_01436_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05928_ (.I(_00899_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05929_ (.I0(\stack[2][3] ),
    .I1(\stack[3][3] ),
    .S(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05930_ (.I0(\stack[0][3] ),
    .I1(\stack[1][3] ),
    .S(_01438_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05931_ (.A1(_00794_),
    .A2(_01473_),
    .B1(_01474_),
    .B2(_01363_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05932_ (.I(_01302_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05933_ (.I0(\stack[4][3] ),
    .I1(\stack[5][3] ),
    .S(_01417_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05934_ (.I0(\stack[6][3] ),
    .I1(\stack[7][3] ),
    .S(_00821_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05935_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_01478_),
    .B2(_01420_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05936_ (.I(_01274_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05937_ (.A1(_01291_),
    .A2(_01475_),
    .B(_01479_),
    .C(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05938_ (.A1(_01471_),
    .A2(_01481_),
    .B(_01446_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05939_ (.I0(\stack[18][4] ),
    .I1(\stack[19][4] ),
    .I2(\stack[16][4] ),
    .I3(\stack[17][4] ),
    .S0(_00856_),
    .S1(_00793_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05940_ (.A1(_01259_),
    .A2(_01483_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05941_ (.I(_01014_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05942_ (.A1(_00900_),
    .A2(\stack[21][4] ),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05943_ (.A1(_01485_),
    .A2(\stack[20][4] ),
    .B(_01303_),
    .C(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05944_ (.A1(_00900_),
    .A2(\stack[23][4] ),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05945_ (.A1(_01485_),
    .A2(\stack[22][4] ),
    .B(_01298_),
    .C(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05946_ (.A1(_01278_),
    .A2(_01484_),
    .A3(_01487_),
    .A4(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05947_ (.I0(\stack[24][4] ),
    .I1(\stack[25][4] ),
    .S(_01391_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05948_ (.I0(\stack[26][4] ),
    .I1(\stack[27][4] ),
    .S(_01369_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05949_ (.A1(_01363_),
    .A2(_01491_),
    .B1(_01492_),
    .B2(_00844_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05950_ (.I0(\stack[28][4] ),
    .I1(\stack[29][4] ),
    .S(_01329_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05951_ (.I0(\stack[30][4] ),
    .I1(\stack[31][4] ),
    .S(_01374_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05952_ (.A1(_01476_),
    .A2(_01494_),
    .B1(_01495_),
    .B2(_01420_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05953_ (.A1(_01342_),
    .A2(_01493_),
    .B(_01496_),
    .C(_01422_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05954_ (.A1(_01490_),
    .A2(_01497_),
    .B(_01424_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05955_ (.A1(_00940_),
    .A2(\stack[5][4] ),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05956_ (.A1(_01485_),
    .A2(\stack[4][4] ),
    .B(_01467_),
    .C(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05957_ (.A1(_00940_),
    .A2(\stack[7][4] ),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05958_ (.A1(_01485_),
    .A2(\stack[6][4] ),
    .B(_01434_),
    .C(_01501_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05959_ (.I0(\stack[2][4] ),
    .I1(\stack[3][4] ),
    .I2(\stack[0][4] ),
    .I3(\stack[1][4] ),
    .S0(_00868_),
    .S1(_00869_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05960_ (.A1(_01398_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05961_ (.A1(_01480_),
    .A2(_01500_),
    .A3(_01502_),
    .A4(_01504_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05962_ (.I0(\stack[10][4] ),
    .I1(\stack[11][4] ),
    .S(_01417_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05963_ (.I0(\stack[8][4] ),
    .I1(\stack[9][4] ),
    .S(_01472_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05964_ (.A1(_01409_),
    .A2(_01506_),
    .B1(_01507_),
    .B2(_01414_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05965_ (.I0(\stack[12][4] ),
    .I1(\stack[13][4] ),
    .S(_01391_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05966_ (.I0(\stack[14][4] ),
    .I1(\stack[15][4] ),
    .S(_01369_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05967_ (.A1(_01390_),
    .A2(_01509_),
    .B1(_01510_),
    .B2(_01394_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05968_ (.A1(_01282_),
    .A2(_01508_),
    .B(_01511_),
    .C(_01307_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05969_ (.A1(_01505_),
    .A2(_01512_),
    .B(_01446_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05970_ (.A1(_01462_),
    .A2(_01482_),
    .A3(_01498_),
    .A4(_01513_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05971_ (.I0(\stack[26][5] ),
    .I1(\stack[27][5] ),
    .S(_01360_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05972_ (.I0(\stack[24][5] ),
    .I1(\stack[25][5] ),
    .S(_01374_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05973_ (.A1(_01426_),
    .A2(_01515_),
    .B1(_01516_),
    .B2(_01430_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05974_ (.I0(\stack[28][5] ),
    .I1(\stack[29][5] ),
    .S(_01438_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05975_ (.I0(\stack[30][5] ),
    .I1(\stack[31][5] ),
    .S(_01371_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05976_ (.A1(_01467_),
    .A2(_01518_),
    .B1(_01519_),
    .B2(_01298_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05977_ (.A1(_01380_),
    .A2(_01517_),
    .B(_01520_),
    .C(_01436_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05978_ (.I0(\stack[18][5] ),
    .I1(\stack[19][5] ),
    .I2(\stack[16][5] ),
    .I3(\stack[17][5] ),
    .S0(_00800_),
    .S1(_00890_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05979_ (.A1(_01398_),
    .A2(_01522_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05980_ (.I0(\stack[20][5] ),
    .I1(\stack[21][5] ),
    .S(_00791_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05981_ (.I0(\stack[22][5] ),
    .I1(\stack[23][5] ),
    .S(_01403_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05982_ (.A1(_01401_),
    .A2(_01524_),
    .B1(_01525_),
    .B2(_01272_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05983_ (.A1(_01355_),
    .A2(_01523_),
    .A3(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05984_ (.A1(_01521_),
    .A2(_01527_),
    .B(_00852_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05985_ (.I0(\stack[2][5] ),
    .I1(\stack[3][5] ),
    .I2(\stack[0][5] ),
    .I3(\stack[1][5] ),
    .S0(_01371_),
    .S1(_00869_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05986_ (.A1(_01259_),
    .A2(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05987_ (.I0(\stack[4][5] ),
    .I1(\stack[5][5] ),
    .S(_01442_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05988_ (.I0(\stack[6][5] ),
    .I1(\stack[7][5] ),
    .S(_01463_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05989_ (.A1(_01390_),
    .A2(_01531_),
    .B1(_01532_),
    .B2(_01394_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05990_ (.A1(_01480_),
    .A2(_01530_),
    .A3(_01533_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05991_ (.I0(\stack[10][5] ),
    .I1(\stack[11][5] ),
    .S(_01463_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05992_ (.I0(\stack[8][5] ),
    .I1(\stack[9][5] ),
    .S(_01427_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05993_ (.A1(_01426_),
    .A2(_01535_),
    .B1(_01536_),
    .B2(_01430_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05994_ (.I0(\stack[12][5] ),
    .I1(\stack[13][5] ),
    .S(_01410_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05995_ (.I0(\stack[14][5] ),
    .I1(\stack[15][5] ),
    .S(_00770_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05996_ (.A1(_01467_),
    .A2(_01538_),
    .B1(_01539_),
    .B2(_01434_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05997_ (.A1(_01380_),
    .A2(_01537_),
    .B(_01540_),
    .C(_01436_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05998_ (.A1(_01534_),
    .A2(_01541_),
    .B(_01446_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05999_ (.I0(\stack[18][1] ),
    .I1(\stack[19][1] ),
    .I2(\stack[16][1] ),
    .I3(\stack[17][1] ),
    .S0(_00827_),
    .S1(_00828_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06000_ (.A1(_01313_),
    .A2(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06001_ (.I0(\stack[22][1] ),
    .I1(\stack[23][1] ),
    .S(_00791_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06002_ (.I0(\stack[20][1] ),
    .I1(\stack[21][1] ),
    .S(_01329_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06003_ (.A1(_01272_),
    .A2(_01545_),
    .B1(_01546_),
    .B2(_01390_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06004_ (.A1(_01275_),
    .A2(_01544_),
    .A3(_01547_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06005_ (.I0(\stack[26][1] ),
    .I1(\stack[27][1] ),
    .S(_01412_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06006_ (.I0(\stack[24][1] ),
    .I1(\stack[25][1] ),
    .S(_01329_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06007_ (.A1(_01409_),
    .A2(_01549_),
    .B1(_01550_),
    .B2(_01414_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06008_ (.I0(\stack[30][1] ),
    .I1(\stack[31][1] ),
    .S(_01391_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06009_ (.I0(\stack[28][1] ),
    .I1(\stack[29][1] ),
    .S(_01438_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06010_ (.A1(_01405_),
    .A2(_01552_),
    .B1(_01553_),
    .B2(_01416_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06011_ (.A1(_01408_),
    .A2(_01551_),
    .B(_01554_),
    .C(_01422_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06012_ (.A1(_01548_),
    .A2(_01555_),
    .B(_01424_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06013_ (.I0(\stack[0][1] ),
    .I1(\stack[1][1] ),
    .S(_01442_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06014_ (.I0(\stack[2][1] ),
    .I1(\stack[3][1] ),
    .S(_01463_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06015_ (.A1(_00931_),
    .A2(_01557_),
    .B1(_01558_),
    .B2(_00891_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06016_ (.I0(\stack[4][1] ),
    .I1(\stack[5][1] ),
    .S(_01472_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06017_ (.I0(\stack[6][1] ),
    .I1(\stack[7][1] ),
    .S(_01374_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06018_ (.A1(_01476_),
    .A2(_01560_),
    .B1(_01561_),
    .B2(_01394_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06019_ (.A1(_01342_),
    .A2(_01559_),
    .B(_01562_),
    .C(_01480_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06020_ (.I0(\stack[10][1] ),
    .I1(\stack[11][1] ),
    .S(_01472_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06021_ (.I0(\stack[8][1] ),
    .I1(\stack[9][1] ),
    .S(_01442_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06022_ (.A1(_01011_),
    .A2(_01564_),
    .B1(_01565_),
    .B2(_01286_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06023_ (.I0(\stack[14][1] ),
    .I1(\stack[15][1] ),
    .S(_00810_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06024_ (.I0(\stack[12][1] ),
    .I1(\stack[13][1] ),
    .S(_01427_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06025_ (.A1(_01405_),
    .A2(_01567_),
    .B1(_01568_),
    .B2(_01476_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06026_ (.A1(_01282_),
    .A2(_01566_),
    .B(_01569_),
    .C(_01307_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06027_ (.A1(_01563_),
    .A2(_01570_),
    .B(_01357_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06028_ (.A1(_01528_),
    .A2(_01542_),
    .A3(_01556_),
    .A4(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06029_ (.A1(_01359_),
    .A2(_01448_),
    .A3(_01514_),
    .A4(_01572_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06030_ (.A1(_01322_),
    .A2(_01573_),
    .B(_01236_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06031_ (.I(_01574_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06032_ (.A1(_01575_),
    .A2(_01232_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06033_ (.A1(_01193_),
    .A2(_01234_),
    .A3(_01219_),
    .A4(_01235_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06034_ (.I(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06035_ (.I(_01322_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06036_ (.A1(_01578_),
    .A2(_01579_),
    .A3(_01573_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06037_ (.A1(_01231_),
    .A2(_01253_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06038_ (.I(_01581_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06039_ (.I(_01252_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06040_ (.A1(_01321_),
    .A2(_01240_),
    .B1(_01583_),
    .B2(_00778_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06041_ (.A1(_01582_),
    .A2(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06042_ (.A1(_01126_),
    .A2(_01576_),
    .B1(_01580_),
    .B2(_01321_),
    .C(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06043_ (.A1(_01254_),
    .A2(_01257_),
    .B(_01586_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06044_ (.I(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06045_ (.A1(_01574_),
    .A2(_01231_),
    .B(_01102_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06046_ (.I(_01239_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06047_ (.A1(_01577_),
    .A2(_01322_),
    .A3(_01573_),
    .B(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06048_ (.A1(_01260_),
    .A2(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06049_ (.A1(_01087_),
    .A2(_01252_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06050_ (.A1(_01581_),
    .A2(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06051_ (.A1(_01036_),
    .A2(_01033_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06052_ (.A1(_01589_),
    .A2(_01592_),
    .A3(_01594_),
    .B1(_01595_),
    .B2(_01581_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06053_ (.I(_01596_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06054_ (.I(_01597_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06055_ (.A1(_01144_),
    .A2(_01591_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06056_ (.A1(_01574_),
    .A2(_01232_),
    .B(_01064_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06057_ (.A1(_01114_),
    .A2(_01583_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06058_ (.A1(_01581_),
    .A2(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06059_ (.A1(_01599_),
    .A2(_01600_),
    .A3(_01602_),
    .B1(_01582_),
    .B2(_01064_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06060_ (.I(_01603_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06061_ (.A1(_01598_),
    .A2(_01604_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06062_ (.I(_01603_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06063_ (.A1(_01597_),
    .A2(_01606_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06064_ (.A1(_01575_),
    .A2(_01232_),
    .B(_01089_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06065_ (.A1(_01279_),
    .A2(_01591_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06066_ (.A1(_01255_),
    .A2(_01583_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06067_ (.A1(_01582_),
    .A2(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06068_ (.A1(_01093_),
    .A2(_01080_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06069_ (.A1(_00805_),
    .A2(_01612_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06070_ (.A1(_01608_),
    .A2(_01609_),
    .A3(_01611_),
    .B1(_01613_),
    .B2(_01582_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06071_ (.I(_01614_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06072_ (.A1(_01607_),
    .A2(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06073_ (.A1(_01588_),
    .A2(_01605_),
    .A3(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06074_ (.I(_01617_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06075_ (.A1(_01583_),
    .A2(_01591_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06076_ (.A1(_01150_),
    .A2(_01619_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06077_ (.A1(_01603_),
    .A2(_01620_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06078_ (.I(net110),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06079_ (.I(net256),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06080_ (.A1(net143),
    .A2(_01623_),
    .A3(net141),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06081_ (.I(net17),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06082_ (.I(net68),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06083_ (.A1(net42),
    .A2(net67),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06084_ (.A1(_01626_),
    .A2(net16),
    .A3(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06085_ (.A1(_01625_),
    .A2(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06086_ (.I(_01629_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06087_ (.A1(_01624_),
    .A2(_01630_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06088_ (.A1(_01622_),
    .A2(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06089_ (.I(_01632_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06090_ (.I(_01251_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06091_ (.I(_01634_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06092_ (.A1(_01633_),
    .A2(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06093_ (.I(_01636_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06094_ (.A1(_01621_),
    .A2(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06095_ (.I(_01638_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06096_ (.I(_01639_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06097_ (.A1(_01618_),
    .A2(_01640_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06098_ (.I(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06099_ (.I(net110),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06100_ (.I(_01643_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06101_ (.A1(_01578_),
    .A2(_01590_),
    .A3(_01204_),
    .A4(_01244_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06102_ (.A1(_01575_),
    .A2(_01645_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06103_ (.A1(_01632_),
    .A2(_01646_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06104_ (.I(_01647_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06105_ (.I(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06106_ (.A1(_01596_),
    .A2(_01603_),
    .A3(_01614_),
    .A4(_01620_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06107_ (.A1(_01587_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06108_ (.A1(_01633_),
    .A2(_01646_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06109_ (.A1(net110),
    .A2(_01629_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06110_ (.I(_01653_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06111_ (.I(net17),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06112_ (.A1(net18),
    .A2(net29),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06113_ (.A1(net1),
    .A2(net2),
    .B(net17),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06114_ (.A1(_01654_),
    .A2(_01655_),
    .B(_01656_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06115_ (.I0(net34),
    .I1(net3),
    .S(net17),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06116_ (.A1(_01657_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06117_ (.I0(net35),
    .I1(net4),
    .S(_01654_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06118_ (.A1(_01659_),
    .A2(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06119_ (.I0(net36),
    .I1(net5),
    .S(_01625_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06120_ (.I0(net38),
    .I1(net7),
    .S(_01654_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06121_ (.I0(net37),
    .I1(net6),
    .S(_01654_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06122_ (.A1(_01663_),
    .A2(_01664_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06123_ (.A1(_01662_),
    .A2(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06124_ (.A1(_01661_),
    .A2(_01666_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06125_ (.A1(prev_reg_write),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06126_ (.A1(_00699_),
    .A2(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06127_ (.I(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06128_ (.I(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06129_ (.A1(_01126_),
    .A2(_01670_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06130_ (.A1(_00850_),
    .A2(_01671_),
    .B(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06131_ (.A1(_01652_),
    .A2(_01673_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06132_ (.A1(_01649_),
    .A2(_01651_),
    .B(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06133_ (.I(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06134_ (.I(_01676_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06135_ (.A1(_01598_),
    .A2(_01621_),
    .B(_01615_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06136_ (.I(_01652_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06137_ (.A1(_01679_),
    .A2(_01650_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06138_ (.A1(_01255_),
    .A2(_01671_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06139_ (.A1(_01137_),
    .A2(_01671_),
    .B(_01681_),
    .C(_01648_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06140_ (.A1(_01678_),
    .A2(_01680_),
    .B(_01682_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06141_ (.I(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06142_ (.I(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06143_ (.A1(_01597_),
    .A2(_01621_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06144_ (.A1(_01127_),
    .A2(_01670_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06145_ (.A1(_01133_),
    .A2(_01671_),
    .B(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06146_ (.I(_01647_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06147_ (.I0(_01686_),
    .I1(_01688_),
    .S(_01689_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06148_ (.I(_01690_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06149_ (.I(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06150_ (.A1(_00699_),
    .A2(_01668_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06151_ (.I(_01666_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06152_ (.I(_01657_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(_01695_),
    .A2(_01658_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06154_ (.A1(_01660_),
    .A2(_01696_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06155_ (.A1(_00699_),
    .A2(_01694_),
    .A3(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06156_ (.A1(_01689_),
    .A2(_01693_),
    .A3(_01698_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06157_ (.I(_01113_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06158_ (.A1(_01700_),
    .A2(_01619_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06159_ (.A1(_01700_),
    .A2(_01670_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06160_ (.I0(_01701_),
    .I1(_01702_),
    .S(_01648_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06161_ (.A1(_01699_),
    .A2(_01703_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06162_ (.A1(_01113_),
    .A2(_01669_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06163_ (.A1(_01130_),
    .A2(_01705_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06164_ (.I(_01620_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06165_ (.A1(_01606_),
    .A2(_01707_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06166_ (.A1(_01606_),
    .A2(_01707_),
    .B(_01647_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06167_ (.A1(_01689_),
    .A2(_01706_),
    .B1(_01708_),
    .B2(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06168_ (.I(_01710_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06169_ (.A1(_01704_),
    .A2(_01711_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06170_ (.I(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06171_ (.A1(_01677_),
    .A2(_01685_),
    .A3(_01692_),
    .A4(_01713_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06172_ (.I(_01638_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06173_ (.A1(_01618_),
    .A2(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06174_ (.A1(_01644_),
    .A2(_01714_),
    .A3(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06175_ (.I(_01717_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06176_ (.I(_01679_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06177_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06178_ (.I(_01625_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06179_ (.I(_01721_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06180_ (.I(_01625_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06181_ (.I(_01723_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06182_ (.I(net8),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06183_ (.A1(_01724_),
    .A2(_01725_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06184_ (.A1(_01722_),
    .A2(net43),
    .B(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06185_ (.I(_01578_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06186_ (.A1(_01728_),
    .A2(_01210_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06187_ (.A1(_01221_),
    .A2(_01729_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06188_ (.I(_01730_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06189_ (.I(_01230_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06190_ (.A1(_01202_),
    .A2(_01245_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06191_ (.A1(_01225_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06192_ (.A1(_01732_),
    .A2(_01634_),
    .A3(_01734_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06193_ (.A1(_01249_),
    .A2(_01731_),
    .A3(_01735_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06194_ (.I(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06195_ (.I(_01359_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06196_ (.A1(_00839_),
    .A2(_01578_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06197_ (.A1(_01738_),
    .A2(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06198_ (.A1(_01738_),
    .A2(_01739_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06199_ (.A1(_01740_),
    .A2(_01741_),
    .B(_01730_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06200_ (.I(_01736_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06201_ (.I(_01246_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06202_ (.I(_01247_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06203_ (.I(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06204_ (.A1(\exec.memory_input[0] ),
    .A2(_01744_),
    .B1(_01746_),
    .B2(_00877_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06205_ (.I(_01635_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06206_ (.A1(_01202_),
    .A2(_01245_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06207_ (.A1(_01732_),
    .A2(_01749_),
    .B(_01181_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06208_ (.A1(_01181_),
    .A2(_01734_),
    .B(_01738_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06209_ (.A1(_01225_),
    .A2(_01748_),
    .A3(_01750_),
    .B(_01751_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06210_ (.A1(_01742_),
    .A2(_01743_),
    .A3(_01747_),
    .A4(_01752_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06211_ (.I(_01719_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06212_ (.A1(_01197_),
    .A2(_01737_),
    .B(_01753_),
    .C(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06213_ (.A1(_01720_),
    .A2(_01727_),
    .B(_01755_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06214_ (.I(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06215_ (.I(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06216_ (.I(_01714_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06217_ (.A1(\stack[2][0] ),
    .A2(_01718_),
    .B1(_01758_),
    .B2(_01759_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06218_ (.A1(_01183_),
    .A2(_01642_),
    .B(_01760_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06219_ (.I(_00874_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06220_ (.I(_01761_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06221_ (.I(_01762_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06222_ (.I(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06223_ (.I(_01721_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06224_ (.I(net9),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06225_ (.I(_01723_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06226_ (.A1(_01766_),
    .A2(_01767_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06227_ (.A1(net54),
    .A2(_01765_),
    .B(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06228_ (.I(_01729_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_01556_),
    .A2(_01571_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06230_ (.I(_01205_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06231_ (.A1(_00838_),
    .A2(_01761_),
    .B(_01236_),
    .C(_01205_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06232_ (.A1(_00840_),
    .A2(_00875_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06233_ (.A1(_00875_),
    .A2(_01772_),
    .B1(_01773_),
    .B2(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06234_ (.A1(_01771_),
    .A2(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06235_ (.A1(_01740_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06236_ (.A1(_01770_),
    .A2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06237_ (.I(_01248_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06238_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06239_ (.A1(\exec.memory_input[1] ),
    .A2(_01744_),
    .B1(_01780_),
    .B2(_00841_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06240_ (.I(_01771_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06241_ (.A1(_00876_),
    .A2(_01782_),
    .A3(_01735_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06242_ (.A1(_01226_),
    .A2(_01634_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06243_ (.A1(_01226_),
    .A2(_01749_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06244_ (.A1(_00876_),
    .A2(_01785_),
    .B(_01782_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06245_ (.A1(_01761_),
    .A2(_01784_),
    .B(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06246_ (.A1(_00918_),
    .A2(_01746_),
    .B1(_01783_),
    .B2(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06247_ (.A1(_01743_),
    .A2(_01781_),
    .A3(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06248_ (.A1(_01211_),
    .A2(_01737_),
    .B1(_01778_),
    .B2(_01789_),
    .C(_01719_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06249_ (.A1(_01720_),
    .A2(_01769_),
    .B(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06250_ (.I(_01791_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06251_ (.I(_01792_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06252_ (.A1(\stack[2][1] ),
    .A2(_01718_),
    .B1(_01793_),
    .B2(_01759_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06253_ (.A1(_01764_),
    .A2(_01642_),
    .B(_01794_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06254_ (.I(_00916_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06255_ (.I(_01795_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06256_ (.I(_01796_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06257_ (.I(net10),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06258_ (.A1(_01724_),
    .A2(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06259_ (.A1(_01722_),
    .A2(net59),
    .B(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06260_ (.I(_01729_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06261_ (.A1(_01782_),
    .A2(_01775_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06262_ (.A1(_01740_),
    .A2(_01776_),
    .B(_01802_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06263_ (.A1(_00917_),
    .A2(_01773_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06264_ (.A1(_01728_),
    .A2(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06265_ (.A1(_01579_),
    .A2(_01805_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06266_ (.A1(_01803_),
    .A2(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06267_ (.I(_01784_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06268_ (.A1(_01732_),
    .A2(_01634_),
    .A3(_01734_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06269_ (.A1(_00916_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06270_ (.I(_01785_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06271_ (.A1(_00918_),
    .A2(_01811_),
    .B(_01579_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06272_ (.A1(_01795_),
    .A2(_01808_),
    .B1(_01810_),
    .B2(_01579_),
    .C(_01812_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06273_ (.I(_00981_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06274_ (.I(_01746_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06275_ (.I(_01736_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06276_ (.A1(\exec.memory_input[2] ),
    .A2(_01744_),
    .B1(_01779_),
    .B2(_00877_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06277_ (.A1(_01814_),
    .A2(_01815_),
    .B(_01816_),
    .C(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06278_ (.A1(_01801_),
    .A2(_01807_),
    .B(_01813_),
    .C(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06279_ (.I(_01736_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06280_ (.I(_01719_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06281_ (.A1(_01228_),
    .A2(_01820_),
    .B(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06282_ (.A1(_01720_),
    .A2(_01800_),
    .B1(_01819_),
    .B2(_01822_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06283_ (.I(_01823_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06284_ (.I(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06285_ (.A1(\stack[2][2] ),
    .A2(_01718_),
    .B1(_01825_),
    .B2(_01759_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06286_ (.A1(_01797_),
    .A2(_01642_),
    .B(_01826_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06287_ (.I(_01814_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06288_ (.I(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06289_ (.I(_01828_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06290_ (.I(_01717_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06291_ (.I(net11),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06292_ (.A1(_01767_),
    .A2(_01831_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06293_ (.A1(_01722_),
    .A2(net60),
    .B(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06294_ (.A1(_01462_),
    .A2(_01482_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06295_ (.I(_01834_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06296_ (.A1(_01357_),
    .A2(_01277_),
    .A3(_01294_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06297_ (.A1(_01357_),
    .A2(_01320_),
    .B(_01836_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06298_ (.A1(_01728_),
    .A2(_01804_),
    .B(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06299_ (.A1(_01803_),
    .A2(_01806_),
    .B(_01838_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06300_ (.A1(_01191_),
    .A2(_01228_),
    .A3(_01237_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06301_ (.A1(_00841_),
    .A2(_00875_),
    .A3(_00917_),
    .B(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06302_ (.I(_01236_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06303_ (.A1(_00981_),
    .A2(_01841_),
    .B(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06304_ (.A1(_00981_),
    .A2(_01841_),
    .B(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06305_ (.A1(_01835_),
    .A2(_01839_),
    .A3(_01844_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06306_ (.I(_01246_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06307_ (.A1(\exec.memory_input[3] ),
    .A2(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06308_ (.A1(_01026_),
    .A2(_01745_),
    .B1(_01779_),
    .B2(_00918_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06309_ (.A1(_01816_),
    .A2(_01847_),
    .A3(_01848_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06310_ (.A1(_01814_),
    .A2(_01809_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06311_ (.A1(_00982_),
    .A2(_01811_),
    .B(_01835_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06312_ (.A1(_01814_),
    .A2(_01808_),
    .B1(_01850_),
    .B2(_01835_),
    .C(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06313_ (.A1(_01801_),
    .A2(_01845_),
    .B(_01849_),
    .C(_01852_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06314_ (.A1(_01191_),
    .A2(_01820_),
    .B(_01754_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06315_ (.A1(_01720_),
    .A2(_01833_),
    .B1(_01853_),
    .B2(_01854_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06316_ (.I(_01855_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06317_ (.I(_01856_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06318_ (.A1(\stack[2][3] ),
    .A2(_01830_),
    .B1(_01857_),
    .B2(_01759_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06319_ (.A1(_01829_),
    .A2(_01642_),
    .B(_01858_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06320_ (.I(_01023_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06321_ (.I(_01859_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06322_ (.I(_01860_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06323_ (.I(net12),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06324_ (.A1(_01721_),
    .A2(_01862_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06325_ (.A1(_01724_),
    .A2(net61),
    .B(_01863_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06326_ (.A1(_01498_),
    .A2(_01513_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06327_ (.I(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06328_ (.A1(_01842_),
    .A2(_01772_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06329_ (.A1(_00839_),
    .A2(_01761_),
    .A3(_00916_),
    .A4(_00980_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06330_ (.A1(_01867_),
    .A2(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06331_ (.A1(_01024_),
    .A2(_01728_),
    .B1(_01867_),
    .B2(_01868_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06332_ (.A1(_01025_),
    .A2(_01869_),
    .B(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06333_ (.A1(_01866_),
    .A2(_01871_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06334_ (.A1(_01834_),
    .A2(_01844_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06335_ (.A1(_01803_),
    .A2(_01806_),
    .B1(_01844_),
    .B2(_01834_),
    .C(_01838_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06336_ (.A1(_01873_),
    .A2(_01874_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06337_ (.A1(_01872_),
    .A2(_01875_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06338_ (.A1(_01026_),
    .A2(_01811_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06339_ (.I(_01866_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06340_ (.A1(_01023_),
    .A2(_01878_),
    .A3(_01809_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06341_ (.A1(_01859_),
    .A2(_01808_),
    .B1(_01877_),
    .B2(_01878_),
    .C(_01879_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(\exec.memory_input[4] ),
    .A2(_01846_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06343_ (.A1(_01074_),
    .A2(_01745_),
    .B1(_01780_),
    .B2(_00983_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06344_ (.A1(_01743_),
    .A2(_01881_),
    .A3(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06345_ (.A1(_01801_),
    .A2(_01876_),
    .B(_01880_),
    .C(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06346_ (.A1(_01215_),
    .A2(_01737_),
    .B(_01754_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06347_ (.A1(_01821_),
    .A2(_01864_),
    .B1(_01884_),
    .B2(_01885_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06348_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06349_ (.I(_01887_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06350_ (.A1(\stack[2][4] ),
    .A2(_01830_),
    .B1(_01888_),
    .B2(_01714_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06351_ (.A1(_01861_),
    .A2(_01641_),
    .B(_01889_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06352_ (.I(_01072_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06353_ (.I(_01890_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06354_ (.I(_01891_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06355_ (.I(_01892_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06356_ (.I(net13),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06357_ (.A1(_01767_),
    .A2(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06358_ (.A1(_01722_),
    .A2(net62),
    .B(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06359_ (.A1(_01865_),
    .A2(_01871_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06360_ (.A1(_01873_),
    .A2(_01897_),
    .A3(_01874_),
    .B1(_01871_),
    .B2(_01866_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06361_ (.A1(_01025_),
    .A2(_01868_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06362_ (.A1(_01772_),
    .A2(_01899_),
    .B(_01890_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06363_ (.I(_01842_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06364_ (.A1(_01072_),
    .A2(_01772_),
    .A3(_01899_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06365_ (.A1(_01901_),
    .A2(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06366_ (.A1(_01528_),
    .A2(_01542_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06367_ (.A1(_01900_),
    .A2(_01903_),
    .B(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06368_ (.A1(_01528_),
    .A2(_01542_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06369_ (.A1(_01025_),
    .A2(_01868_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06370_ (.A1(_01840_),
    .A2(_01907_),
    .B(_01073_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06371_ (.A1(_01842_),
    .A2(_01906_),
    .A3(_01908_),
    .A4(_01902_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06372_ (.I(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06373_ (.A1(_01905_),
    .A2(_01910_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06374_ (.A1(_01898_),
    .A2(_01911_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06375_ (.A1(\exec.memory_input[5] ),
    .A2(_01744_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06376_ (.A1(_01122_),
    .A2(_01745_),
    .B1(_01779_),
    .B2(_01026_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06377_ (.A1(_01816_),
    .A2(_01913_),
    .A3(_01914_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06378_ (.A1(_01074_),
    .A2(_01811_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06379_ (.A1(_01890_),
    .A2(_01904_),
    .A3(_01809_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06380_ (.A1(_01890_),
    .A2(_01808_),
    .B1(_01916_),
    .B2(_01904_),
    .C(_01917_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06381_ (.A1(_01729_),
    .A2(_01912_),
    .B(_01915_),
    .C(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06382_ (.A1(_01233_),
    .A2(_01737_),
    .B(_01754_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06383_ (.A1(_01821_),
    .A2(_01896_),
    .B1(_01919_),
    .B2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06384_ (.I(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06385_ (.I(_01922_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06386_ (.A1(\stack[2][5] ),
    .A2(_01830_),
    .B1(_01923_),
    .B2(_01714_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06387_ (.A1(_01893_),
    .A2(_01641_),
    .B(_01924_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06388_ (.I(_01684_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06389_ (.A1(_01677_),
    .A2(_01925_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06390_ (.A1(_01648_),
    .A2(_01688_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06391_ (.A1(_01679_),
    .A2(_01686_),
    .B(_01927_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06392_ (.I(_01928_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06393_ (.I(_01929_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06394_ (.I(_01930_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06395_ (.A1(_01926_),
    .A2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06396_ (.I(_01713_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06397_ (.A1(_01932_),
    .A2(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06398_ (.A1(_01425_),
    .A2(_01447_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06399_ (.I(_01121_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06400_ (.I(_01936_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06401_ (.A1(_01073_),
    .A2(_01907_),
    .B(_01840_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06402_ (.A1(_01936_),
    .A2(_01938_),
    .B(_01901_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06403_ (.A1(_01937_),
    .A2(_01938_),
    .B(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06404_ (.A1(_01935_),
    .A2(_01940_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06405_ (.A1(_01901_),
    .A2(_01908_),
    .A3(_01902_),
    .B(_01906_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06406_ (.A1(_01872_),
    .A2(_01942_),
    .A3(_01909_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _06407_ (.A1(_01878_),
    .A2(_01871_),
    .A3(_01910_),
    .B1(_01943_),
    .B2(_01874_),
    .B3(_01873_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06408_ (.A1(_01905_),
    .A2(_01941_),
    .A3(_01944_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06409_ (.A1(_01905_),
    .A2(_01944_),
    .B(_01941_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06410_ (.A1(_01801_),
    .A2(_01945_),
    .A3(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06411_ (.A1(\exec.memory_input[6] ),
    .A2(_01846_),
    .B1(_01746_),
    .B2(_01169_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06412_ (.I(_01935_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06413_ (.A1(_01123_),
    .A2(_01949_),
    .A3(_01735_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06414_ (.A1(_01122_),
    .A2(_01785_),
    .B(_01949_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06415_ (.A1(_01937_),
    .A2(_01784_),
    .B(_01951_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06416_ (.A1(_01075_),
    .A2(_01780_),
    .B1(_01950_),
    .B2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06417_ (.A1(_01743_),
    .A2(_01948_),
    .A3(_01953_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06418_ (.A1(_01217_),
    .A2(_01820_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06419_ (.A1(_01947_),
    .A2(_01954_),
    .B(_01955_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06420_ (.I(net14),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06421_ (.A1(_01723_),
    .A2(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06422_ (.A1(_01721_),
    .A2(net63),
    .B(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06423_ (.I(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06424_ (.A1(_01649_),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06425_ (.A1(_01649_),
    .A2(_01956_),
    .B(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06426_ (.I(_01962_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06427_ (.I(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06428_ (.A1(\stack[2][6] ),
    .A2(_01718_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06429_ (.A1(net151),
    .A2(_01716_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06430_ (.A1(_01934_),
    .A2(_01964_),
    .B(_01965_),
    .C(_01966_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(_01949_),
    .A2(_01940_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06432_ (.A1(_01379_),
    .A2(_01397_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06433_ (.A1(_01074_),
    .A2(_01122_),
    .A3(_01907_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06434_ (.A1(_01168_),
    .A2(_01901_),
    .B1(_01867_),
    .B2(_01969_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06435_ (.A1(_01167_),
    .A2(_01968_),
    .A3(_01970_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06436_ (.A1(_01967_),
    .A2(_01946_),
    .A3(_01971_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06437_ (.A1(_01967_),
    .A2(_01946_),
    .B(_01971_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06438_ (.I(_01780_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06439_ (.I(_01167_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06440_ (.A1(_01937_),
    .A2(_01974_),
    .B1(_01749_),
    .B2(_01975_),
    .C(_01816_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06441_ (.A1(_01168_),
    .A2(_01968_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06442_ (.A1(_01379_),
    .A2(_01397_),
    .B(_01225_),
    .C(_01975_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06443_ (.A1(_01975_),
    .A2(_01732_),
    .B(_01635_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06444_ (.A1(_01968_),
    .A2(_01979_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06445_ (.A1(_01226_),
    .A2(_01977_),
    .A3(_01978_),
    .B(_01980_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06446_ (.A1(\exec.memory_input[7] ),
    .A2(_01846_),
    .B(_01976_),
    .C(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06447_ (.A1(_01770_),
    .A2(_01972_),
    .A3(_01973_),
    .B(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06448_ (.A1(_01216_),
    .A2(_01820_),
    .B(_01821_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06449_ (.I(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06450_ (.I(net15),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06451_ (.A1(_01765_),
    .A2(net64),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06452_ (.A1(_01765_),
    .A2(_01986_),
    .B(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06453_ (.A1(_01983_),
    .A2(_01985_),
    .B1(_01988_),
    .B2(_01649_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06454_ (.I(_01989_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06455_ (.I(_01990_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06456_ (.A1(net152),
    .A2(_01716_),
    .B1(_01830_),
    .B2(\stack[2][7] ),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06457_ (.A1(_01934_),
    .A2(_01991_),
    .B(_01992_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06458_ (.I(_01177_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06459_ (.A1(_00763_),
    .A2(_01172_),
    .A3(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06460_ (.I(_01994_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06461_ (.A1(\mem.mem_dff.cycles[1] ),
    .A2(\mem.mem_dff.cycles[0] ),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06462_ (.I(_01622_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06463_ (.I(_01997_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06464_ (.I(_01998_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06465_ (.I(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06466_ (.A1(\mem.dff_data_ready ),
    .A2(_01996_),
    .B(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06467_ (.A1(_01995_),
    .A2(_02001_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06468_ (.I(_01643_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06469_ (.I(_02002_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06470_ (.I(_02003_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06471_ (.I(_02004_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06472_ (.A1(\mem.mem_dff.cycles[0] ),
    .A2(_01995_),
    .A3(_01996_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06473_ (.A1(\mem.mem_dff.cycles[0] ),
    .A2(_01995_),
    .B(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06474_ (.A1(_02005_),
    .A2(_02007_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06475_ (.I(_01997_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06476_ (.I(_02008_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06477_ (.I(_02009_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06478_ (.A1(\mem.mem_dff.cycles[1] ),
    .A2(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06479_ (.A1(_02006_),
    .A2(_02011_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06480_ (.I(\mem.mem_dff.code_mem[0][0] ),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06481_ (.A1(net253),
    .A2(_01996_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06482_ (.A1(_01994_),
    .A2(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06483_ (.A1(_00764_),
    .A2(_01175_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06484_ (.A1(_02014_),
    .A2(_02015_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06485_ (.I(_02016_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06486_ (.I(_02017_),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06487_ (.I(net255),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06488_ (.I(_02019_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06489_ (.A1(_02020_),
    .A2(net227),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06490_ (.I(net187),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06491_ (.I(net254),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06492_ (.A1(_02022_),
    .A2(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06493_ (.I(_02024_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06494_ (.A1(_02021_),
    .A2(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06495_ (.I(_02026_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06496_ (.A1(_02018_),
    .A2(_02027_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06497_ (.I(_02028_),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06498_ (.I(net249),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06499_ (.I(_02030_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06500_ (.I(_02028_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06501_ (.I(_01999_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06502_ (.A1(_02031_),
    .A2(_02032_),
    .B(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06503_ (.A1(_02012_),
    .A2(_02029_),
    .B(_02034_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06504_ (.I(\mem.mem_dff.code_mem[0][1] ),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06505_ (.I(net248),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06506_ (.I(_02036_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06507_ (.A1(_02037_),
    .A2(_02032_),
    .B(_02033_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06508_ (.A1(_02035_),
    .A2(_02029_),
    .B(_02038_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06509_ (.I(\mem.mem_dff.code_mem[0][2] ),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06510_ (.I(net244),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06511_ (.I(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06512_ (.A1(_02041_),
    .A2(_02032_),
    .B(_02033_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06513_ (.A1(_02039_),
    .A2(_02029_),
    .B(_02042_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06514_ (.I(\mem.mem_dff.code_mem[0][3] ),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06515_ (.I(net242),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06516_ (.I(_02044_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06517_ (.I(_01999_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06518_ (.A1(_02045_),
    .A2(_02032_),
    .B(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06519_ (.A1(_02043_),
    .A2(_02029_),
    .B(_02047_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06520_ (.I(\mem.mem_dff.code_mem[0][4] ),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06521_ (.I(_02028_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06522_ (.I(net241),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06523_ (.I(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06524_ (.I(_02028_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06525_ (.A1(_02051_),
    .A2(_02052_),
    .B(_02046_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06526_ (.A1(_02048_),
    .A2(_02049_),
    .B(_02053_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06527_ (.I(\mem.mem_dff.code_mem[0][5] ),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06528_ (.I(net237),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06529_ (.I(_02055_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06530_ (.A1(_02056_),
    .A2(_02052_),
    .B(_02046_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06531_ (.A1(_02054_),
    .A2(_02049_),
    .B(_02057_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06532_ (.I(\mem.mem_dff.code_mem[0][6] ),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06533_ (.I(net235),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06534_ (.I(_02059_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06535_ (.A1(_02060_),
    .A2(_02052_),
    .B(_02046_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06536_ (.A1(_02058_),
    .A2(_02049_),
    .B(_02061_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06537_ (.I(\mem.mem_dff.code_mem[0][7] ),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06538_ (.I(net233),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06539_ (.I(_02063_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06540_ (.I(_02008_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06541_ (.I(_02065_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06542_ (.A1(_02064_),
    .A2(_02052_),
    .B(_02066_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06543_ (.A1(_02062_),
    .A2(_02049_),
    .B(_02067_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06544_ (.I(\mem.mem_dff.code_mem[1][0] ),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06545_ (.A1(_02019_),
    .A2(net228),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06546_ (.A1(_02025_),
    .A2(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06547_ (.I(_02070_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06548_ (.A1(_02018_),
    .A2(_02071_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06549_ (.I(_02072_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06550_ (.I(_02072_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06551_ (.A1(_02031_),
    .A2(_02074_),
    .B(_02066_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06552_ (.A1(_02068_),
    .A2(_02073_),
    .B(_02075_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06553_ (.I(\mem.mem_dff.code_mem[1][1] ),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06554_ (.A1(_02037_),
    .A2(_02074_),
    .B(_02066_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06555_ (.A1(_02076_),
    .A2(_02073_),
    .B(_02077_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06556_ (.I(\mem.mem_dff.code_mem[1][2] ),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06557_ (.A1(_02041_),
    .A2(_02074_),
    .B(_02066_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06558_ (.A1(_02078_),
    .A2(_02073_),
    .B(_02079_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06559_ (.I(\mem.mem_dff.code_mem[1][3] ),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06560_ (.I(_02065_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06561_ (.A1(_02045_),
    .A2(_02074_),
    .B(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06562_ (.A1(_02080_),
    .A2(_02073_),
    .B(_02082_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06563_ (.I(\mem.mem_dff.code_mem[1][4] ),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06564_ (.I(_02072_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06565_ (.I(_02072_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06566_ (.A1(_02051_),
    .A2(_02085_),
    .B(_02081_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06567_ (.A1(_02083_),
    .A2(_02084_),
    .B(_02086_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06568_ (.I(\mem.mem_dff.code_mem[1][5] ),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06569_ (.A1(_02056_),
    .A2(_02085_),
    .B(_02081_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06570_ (.A1(_02087_),
    .A2(_02084_),
    .B(_02088_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06571_ (.I(\mem.mem_dff.code_mem[1][6] ),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06572_ (.A1(_02060_),
    .A2(_02085_),
    .B(_02081_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06573_ (.A1(_02089_),
    .A2(_02084_),
    .B(_02090_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06574_ (.I(\mem.mem_dff.code_mem[1][7] ),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06575_ (.I(_02065_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06576_ (.A1(_02064_),
    .A2(_02085_),
    .B(_02092_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06577_ (.A1(_02091_),
    .A2(_02084_),
    .B(_02093_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06578_ (.I(\mem.mem_dff.code_mem[2][0] ),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06579_ (.I(_02024_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06580_ (.A1(_02020_),
    .A2(net229),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06581_ (.A1(_02095_),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06582_ (.I(_02097_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06583_ (.A1(_02018_),
    .A2(_02098_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06584_ (.I(_02099_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06585_ (.I(net249),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06586_ (.I(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06587_ (.I(_02099_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06588_ (.A1(_02102_),
    .A2(_02103_),
    .B(_02092_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06589_ (.A1(_02094_),
    .A2(_02100_),
    .B(_02104_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06590_ (.I(\mem.mem_dff.code_mem[2][1] ),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06591_ (.A1(_02037_),
    .A2(_02103_),
    .B(_02092_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06592_ (.A1(_02105_),
    .A2(_02100_),
    .B(_02106_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06593_ (.I(\mem.mem_dff.code_mem[2][2] ),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06594_ (.I(net244),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06595_ (.I(_02108_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06596_ (.A1(_02109_),
    .A2(_02103_),
    .B(_02092_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06597_ (.A1(_02107_),
    .A2(_02100_),
    .B(_02110_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06598_ (.I(\mem.mem_dff.code_mem[2][3] ),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06599_ (.I(_02065_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06600_ (.A1(_02045_),
    .A2(_02103_),
    .B(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06601_ (.A1(_02111_),
    .A2(_02100_),
    .B(_02113_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06602_ (.I(\mem.mem_dff.code_mem[2][4] ),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06603_ (.I(_02099_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06604_ (.I(net240),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06605_ (.I(_02116_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06606_ (.I(_02099_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06607_ (.A1(_02117_),
    .A2(_02118_),
    .B(_02112_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06608_ (.A1(_02114_),
    .A2(_02115_),
    .B(_02119_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06609_ (.I(\mem.mem_dff.code_mem[2][5] ),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06610_ (.I(net237),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06611_ (.I(_02121_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06612_ (.A1(_02122_),
    .A2(_02118_),
    .B(_02112_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06613_ (.A1(_02120_),
    .A2(_02115_),
    .B(_02123_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06614_ (.I(\mem.mem_dff.code_mem[2][6] ),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06615_ (.A1(_02060_),
    .A2(_02118_),
    .B(_02112_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06616_ (.A1(_02124_),
    .A2(_02115_),
    .B(_02125_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06617_ (.I(\mem.mem_dff.code_mem[2][7] ),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06618_ (.I(_01997_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06619_ (.I(_02127_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06620_ (.I(_02128_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06621_ (.I(_02129_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06622_ (.A1(_02064_),
    .A2(_02118_),
    .B(_02130_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06623_ (.A1(_02126_),
    .A2(_02115_),
    .B(_02131_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06624_ (.I(\mem.mem_dff.code_mem[3][0] ),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06625_ (.I(net255),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06626_ (.I(_00759_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06627_ (.I(_02134_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06628_ (.A1(_02133_),
    .A2(_02135_),
    .A3(_02095_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06629_ (.I(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06630_ (.A1(_02018_),
    .A2(_02137_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06631_ (.I(_02138_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06632_ (.I(_02138_),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06633_ (.A1(_02102_),
    .A2(_02140_),
    .B(_02130_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06634_ (.A1(_02132_),
    .A2(_02139_),
    .B(_02141_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06635_ (.I(\mem.mem_dff.code_mem[3][1] ),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06636_ (.I(net247),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06637_ (.I(_02143_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06638_ (.A1(_02144_),
    .A2(_02140_),
    .B(_02130_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06639_ (.A1(_02142_),
    .A2(_02139_),
    .B(_02145_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06640_ (.I(\mem.mem_dff.code_mem[3][2] ),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06641_ (.A1(_02109_),
    .A2(_02140_),
    .B(_02130_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06642_ (.A1(_02146_),
    .A2(_02139_),
    .B(_02147_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06643_ (.I(\mem.mem_dff.code_mem[3][3] ),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06644_ (.I(net242),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06645_ (.I(_02149_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06646_ (.I(_02129_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06647_ (.A1(_02150_),
    .A2(_02140_),
    .B(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06648_ (.A1(_02148_),
    .A2(_02139_),
    .B(_02152_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06649_ (.I(\mem.mem_dff.code_mem[3][4] ),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06650_ (.I(_02138_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06651_ (.I(_02138_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06652_ (.A1(_02117_),
    .A2(_02155_),
    .B(_02151_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06653_ (.A1(_02153_),
    .A2(_02154_),
    .B(_02156_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06654_ (.I(\mem.mem_dff.code_mem[3][5] ),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06655_ (.A1(_02122_),
    .A2(_02155_),
    .B(_02151_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06656_ (.A1(_02157_),
    .A2(_02154_),
    .B(_02158_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06657_ (.I(\mem.mem_dff.code_mem[3][6] ),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(net235),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06659_ (.I(_02160_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06660_ (.A1(_02161_),
    .A2(_02155_),
    .B(_02151_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06661_ (.A1(_02159_),
    .A2(_02154_),
    .B(_02162_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06662_ (.I(\mem.mem_dff.code_mem[3][7] ),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06663_ (.I(net233),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06664_ (.I(_02164_),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06665_ (.I(_02129_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06666_ (.A1(_02165_),
    .A2(_02155_),
    .B(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06667_ (.A1(_02163_),
    .A2(_02154_),
    .B(_02167_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06668_ (.I(\mem.mem_dff.code_mem[4][0] ),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06669_ (.I(_02017_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06670_ (.I(net255),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06671_ (.A1(_02170_),
    .A2(net227),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06672_ (.A1(_02095_),
    .A2(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06673_ (.I(_02172_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06674_ (.A1(_02169_),
    .A2(_02173_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06675_ (.I(_02174_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06676_ (.I(_02174_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06677_ (.A1(_02102_),
    .A2(_02176_),
    .B(_02166_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06678_ (.A1(_02168_),
    .A2(_02175_),
    .B(_02177_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06679_ (.I(\mem.mem_dff.code_mem[4][1] ),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06680_ (.A1(_02144_),
    .A2(_02176_),
    .B(_02166_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06681_ (.A1(_02178_),
    .A2(_02175_),
    .B(_02179_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06682_ (.I(\mem.mem_dff.code_mem[4][2] ),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06683_ (.A1(_02109_),
    .A2(_02176_),
    .B(_02166_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06684_ (.A1(_02180_),
    .A2(_02175_),
    .B(_02181_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06685_ (.I(\mem.mem_dff.code_mem[4][3] ),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06686_ (.I(_02129_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06687_ (.A1(_02150_),
    .A2(_02176_),
    .B(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06688_ (.A1(_02182_),
    .A2(_02175_),
    .B(_02184_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06689_ (.I(\mem.mem_dff.code_mem[4][4] ),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06690_ (.I(_02174_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06691_ (.I(_02174_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06692_ (.A1(_02117_),
    .A2(_02187_),
    .B(_02183_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06693_ (.A1(_02185_),
    .A2(_02186_),
    .B(_02188_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06694_ (.I(\mem.mem_dff.code_mem[4][5] ),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06695_ (.A1(_02122_),
    .A2(_02187_),
    .B(_02183_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06696_ (.A1(_02189_),
    .A2(_02186_),
    .B(_02190_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06697_ (.I(\mem.mem_dff.code_mem[4][6] ),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06698_ (.A1(_02161_),
    .A2(_02187_),
    .B(_02183_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06699_ (.A1(_02191_),
    .A2(_02186_),
    .B(_02192_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06700_ (.I(\mem.mem_dff.code_mem[4][7] ),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06701_ (.I(_02128_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06702_ (.I(_02194_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06703_ (.A1(_02165_),
    .A2(_02187_),
    .B(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06704_ (.A1(_02193_),
    .A2(_02186_),
    .B(_02196_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06705_ (.I(\mem.mem_dff.code_mem[5][0] ),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06706_ (.A1(_02170_),
    .A2(net228),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06707_ (.A1(_02025_),
    .A2(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06708_ (.I(_02199_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(_02169_),
    .A2(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06710_ (.I(_02201_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06711_ (.I(_02201_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06712_ (.A1(_02102_),
    .A2(_02203_),
    .B(_02195_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06713_ (.A1(_02197_),
    .A2(_02202_),
    .B(_02204_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06714_ (.I(\mem.mem_dff.code_mem[5][1] ),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06715_ (.A1(_02144_),
    .A2(_02203_),
    .B(_02195_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06716_ (.A1(_02205_),
    .A2(_02202_),
    .B(_02206_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06717_ (.I(\mem.mem_dff.code_mem[5][2] ),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06718_ (.A1(_02109_),
    .A2(_02203_),
    .B(_02195_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06719_ (.A1(_02207_),
    .A2(_02202_),
    .B(_02208_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06720_ (.I(\mem.mem_dff.code_mem[5][3] ),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06721_ (.I(_02194_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06722_ (.A1(_02150_),
    .A2(_02203_),
    .B(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06723_ (.A1(_02209_),
    .A2(_02202_),
    .B(_02211_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06724_ (.I(\mem.mem_dff.code_mem[5][4] ),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06725_ (.I(_02201_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06726_ (.I(_02201_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06727_ (.A1(_02117_),
    .A2(_02214_),
    .B(_02210_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06728_ (.A1(_02212_),
    .A2(_02213_),
    .B(_02215_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06729_ (.I(\mem.mem_dff.code_mem[5][5] ),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06730_ (.A1(_02122_),
    .A2(_02214_),
    .B(_02210_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06731_ (.A1(_02216_),
    .A2(_02213_),
    .B(_02217_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06732_ (.I(\mem.mem_dff.code_mem[5][6] ),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06733_ (.A1(_02161_),
    .A2(_02214_),
    .B(_02210_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06734_ (.A1(_02218_),
    .A2(_02213_),
    .B(_02219_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06735_ (.I(\mem.mem_dff.code_mem[5][7] ),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06736_ (.I(_02194_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06737_ (.A1(_02165_),
    .A2(_02214_),
    .B(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06738_ (.A1(_02220_),
    .A2(_02213_),
    .B(_02222_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06739_ (.I(\mem.mem_dff.code_mem[6][0] ),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06740_ (.A1(_02170_),
    .A2(net229),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06741_ (.A1(_02095_),
    .A2(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06742_ (.I(_02225_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_02169_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06744_ (.I(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06745_ (.I(_02101_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06746_ (.I(_02227_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06747_ (.A1(_02229_),
    .A2(_02230_),
    .B(_02221_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06748_ (.A1(_02223_),
    .A2(_02228_),
    .B(_02231_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06749_ (.I(\mem.mem_dff.code_mem[6][1] ),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06750_ (.A1(_02144_),
    .A2(_02230_),
    .B(_02221_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06751_ (.A1(_02232_),
    .A2(_02228_),
    .B(_02233_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06752_ (.I(\mem.mem_dff.code_mem[6][2] ),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06753_ (.I(_02108_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06754_ (.A1(_02235_),
    .A2(_02230_),
    .B(_02221_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06755_ (.A1(_02234_),
    .A2(_02228_),
    .B(_02236_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06756_ (.I(\mem.mem_dff.code_mem[6][3] ),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06757_ (.I(_02194_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06758_ (.A1(_02150_),
    .A2(_02230_),
    .B(_02238_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06759_ (.A1(_02237_),
    .A2(_02228_),
    .B(_02239_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06760_ (.I(\mem.mem_dff.code_mem[6][4] ),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06761_ (.I(_02227_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06762_ (.I(_02116_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06763_ (.I(_02227_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06764_ (.A1(_02242_),
    .A2(_02243_),
    .B(_02238_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06765_ (.A1(_02240_),
    .A2(_02241_),
    .B(_02244_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06766_ (.I(\mem.mem_dff.code_mem[6][5] ),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06767_ (.I(_02121_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06768_ (.A1(_02246_),
    .A2(_02243_),
    .B(_02238_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06769_ (.A1(_02245_),
    .A2(_02241_),
    .B(_02247_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06770_ (.I(\mem.mem_dff.code_mem[6][6] ),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06771_ (.A1(_02161_),
    .A2(_02243_),
    .B(_02238_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06772_ (.A1(_02248_),
    .A2(_02241_),
    .B(_02249_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06773_ (.I(\mem.mem_dff.code_mem[6][7] ),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06774_ (.I(_02128_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06775_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06776_ (.A1(_02165_),
    .A2(_02243_),
    .B(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06777_ (.A1(_02250_),
    .A2(_02241_),
    .B(_02253_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06778_ (.I(\mem.mem_dff.code_mem[7][0] ),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06779_ (.A1(_02170_),
    .A2(net230),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06780_ (.I(_02255_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06781_ (.A1(_02025_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06782_ (.I(_02257_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06783_ (.A1(_02169_),
    .A2(_02258_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06784_ (.I(_02259_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06785_ (.I(_02259_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06786_ (.A1(_02229_),
    .A2(_02261_),
    .B(_02252_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06787_ (.A1(_02254_),
    .A2(_02260_),
    .B(_02262_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06788_ (.I(\mem.mem_dff.code_mem[7][1] ),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06789_ (.I(_02143_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06790_ (.A1(_02264_),
    .A2(_02261_),
    .B(_02252_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06791_ (.A1(_02263_),
    .A2(_02260_),
    .B(_02265_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06792_ (.I(\mem.mem_dff.code_mem[7][2] ),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06793_ (.A1(_02235_),
    .A2(_02261_),
    .B(_02252_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06794_ (.A1(_02266_),
    .A2(_02260_),
    .B(_02267_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06795_ (.I(\mem.mem_dff.code_mem[7][3] ),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06796_ (.I(_02149_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06797_ (.I(_02251_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06798_ (.A1(_02269_),
    .A2(_02261_),
    .B(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06799_ (.A1(_02268_),
    .A2(_02260_),
    .B(_02271_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06800_ (.I(\mem.mem_dff.code_mem[7][4] ),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06801_ (.I(_02259_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06802_ (.I(_02259_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06803_ (.A1(_02242_),
    .A2(_02274_),
    .B(_02270_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06804_ (.A1(_02272_),
    .A2(_02273_),
    .B(_02275_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06805_ (.I(\mem.mem_dff.code_mem[7][5] ),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06806_ (.A1(_02246_),
    .A2(_02274_),
    .B(_02270_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06807_ (.A1(_02276_),
    .A2(_02273_),
    .B(_02277_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06808_ (.I(\mem.mem_dff.code_mem[7][6] ),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06809_ (.I(_02160_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06810_ (.A1(_02279_),
    .A2(_02274_),
    .B(_02270_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06811_ (.A1(_02278_),
    .A2(_02273_),
    .B(_02280_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06812_ (.I(\mem.mem_dff.code_mem[7][7] ),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06813_ (.I(_02164_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06814_ (.I(_02251_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06815_ (.A1(_02282_),
    .A2(_02274_),
    .B(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06816_ (.A1(_02281_),
    .A2(_02273_),
    .B(_02284_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06817_ (.I(\mem.mem_dff.code_mem[8][0] ),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06818_ (.I(_02017_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06819_ (.I(net187),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06820_ (.I(_02287_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06821_ (.I(_00758_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06822_ (.A1(net255),
    .A2(_02289_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(net254),
    .A2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06824_ (.A1(_02288_),
    .A2(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06825_ (.I(_02292_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06826_ (.A1(_02286_),
    .A2(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06827_ (.I(_02294_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06828_ (.I(_02294_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06829_ (.A1(_02229_),
    .A2(_02296_),
    .B(_02283_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06830_ (.A1(_02285_),
    .A2(_02295_),
    .B(_02297_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06831_ (.I(\mem.mem_dff.code_mem[8][1] ),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06832_ (.A1(_02264_),
    .A2(_02296_),
    .B(_02283_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06833_ (.A1(_02298_),
    .A2(_02295_),
    .B(_02299_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06834_ (.I(\mem.mem_dff.code_mem[8][2] ),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06835_ (.A1(_02235_),
    .A2(_02296_),
    .B(_02283_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06836_ (.A1(_02300_),
    .A2(_02295_),
    .B(_02301_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06837_ (.I(\mem.mem_dff.code_mem[8][3] ),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06838_ (.I(_02251_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06839_ (.A1(_02269_),
    .A2(_02296_),
    .B(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06840_ (.A1(_02302_),
    .A2(_02295_),
    .B(_02304_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06841_ (.I(\mem.mem_dff.code_mem[8][4] ),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06842_ (.I(_02294_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06843_ (.I(_02294_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06844_ (.A1(_02242_),
    .A2(_02307_),
    .B(_02303_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06845_ (.A1(_02305_),
    .A2(_02306_),
    .B(_02308_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06846_ (.I(\mem.mem_dff.code_mem[8][5] ),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06847_ (.A1(_02246_),
    .A2(_02307_),
    .B(_02303_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06848_ (.A1(_02309_),
    .A2(_02306_),
    .B(_02310_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06849_ (.I(\mem.mem_dff.code_mem[8][6] ),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06850_ (.A1(_02279_),
    .A2(_02307_),
    .B(_02303_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06851_ (.A1(_02311_),
    .A2(_02306_),
    .B(_02312_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06852_ (.I(\mem.mem_dff.code_mem[8][7] ),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06853_ (.I(_02128_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06854_ (.I(_02314_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06855_ (.A1(_02282_),
    .A2(_02307_),
    .B(_02315_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06856_ (.A1(_02313_),
    .A2(_02306_),
    .B(_02316_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06857_ (.I(\mem.mem_dff.code_mem[9][0] ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06858_ (.I(_02023_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06859_ (.I(_02318_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06860_ (.A1(_02288_),
    .A2(_02319_),
    .A3(_02069_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06861_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06862_ (.A1(_02286_),
    .A2(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06863_ (.I(_02322_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06864_ (.I(_02322_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06865_ (.A1(_02229_),
    .A2(_02324_),
    .B(_02315_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06866_ (.A1(_02317_),
    .A2(_02323_),
    .B(_02325_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06867_ (.I(\mem.mem_dff.code_mem[9][1] ),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06868_ (.A1(_02264_),
    .A2(_02324_),
    .B(_02315_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06869_ (.A1(_02326_),
    .A2(_02323_),
    .B(_02327_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06870_ (.I(\mem.mem_dff.code_mem[9][2] ),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06871_ (.A1(_02235_),
    .A2(_02324_),
    .B(_02315_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06872_ (.A1(_02328_),
    .A2(_02323_),
    .B(_02329_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06873_ (.I(\mem.mem_dff.code_mem[9][3] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06874_ (.I(_02314_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06875_ (.A1(_02269_),
    .A2(_02324_),
    .B(_02331_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06876_ (.A1(_02330_),
    .A2(_02323_),
    .B(_02332_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06877_ (.I(\mem.mem_dff.code_mem[9][4] ),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06878_ (.I(_02322_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06879_ (.I(_02322_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06880_ (.A1(_02242_),
    .A2(_02335_),
    .B(_02331_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06881_ (.A1(_02333_),
    .A2(_02334_),
    .B(_02336_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06882_ (.I(\mem.mem_dff.code_mem[9][5] ),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06883_ (.A1(_02246_),
    .A2(_02335_),
    .B(_02331_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06884_ (.A1(_02337_),
    .A2(_02334_),
    .B(_02338_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06885_ (.I(\mem.mem_dff.code_mem[9][6] ),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06886_ (.A1(_02279_),
    .A2(_02335_),
    .B(_02331_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06887_ (.A1(_02339_),
    .A2(_02334_),
    .B(_02340_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06888_ (.I(\mem.mem_dff.code_mem[9][7] ),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06889_ (.I(_02314_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06890_ (.A1(_02282_),
    .A2(_02335_),
    .B(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06891_ (.A1(_02341_),
    .A2(_02334_),
    .B(_02343_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06892_ (.I(\mem.mem_dff.code_mem[10][0] ),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06893_ (.I(_02287_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06894_ (.A1(_02345_),
    .A2(_02319_),
    .A3(_02096_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06895_ (.I(_02346_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06896_ (.A1(_02286_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06897_ (.I(_02348_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06898_ (.I(net249),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06899_ (.I(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06900_ (.I(_02348_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06901_ (.A1(_02351_),
    .A2(_02352_),
    .B(_02342_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06902_ (.A1(_02344_),
    .A2(_02349_),
    .B(_02353_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06903_ (.I(\mem.mem_dff.code_mem[10][1] ),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06904_ (.A1(_02264_),
    .A2(_02352_),
    .B(_02342_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06905_ (.A1(_02354_),
    .A2(_02349_),
    .B(_02355_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06906_ (.I(\mem.mem_dff.code_mem[10][2] ),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06907_ (.I(net244),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06908_ (.I(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06909_ (.A1(_02358_),
    .A2(_02352_),
    .B(_02342_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06910_ (.A1(_02356_),
    .A2(_02349_),
    .B(_02359_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06911_ (.I(\mem.mem_dff.code_mem[10][3] ),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06912_ (.I(_02314_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06913_ (.A1(_02269_),
    .A2(_02352_),
    .B(_02361_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06914_ (.A1(_02360_),
    .A2(_02349_),
    .B(_02362_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06915_ (.I(\mem.mem_dff.code_mem[10][4] ),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06916_ (.I(_02348_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06917_ (.I(net240),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06918_ (.I(_02365_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06919_ (.I(_02348_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06920_ (.A1(_02366_),
    .A2(_02367_),
    .B(_02361_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06921_ (.A1(_02363_),
    .A2(_02364_),
    .B(_02368_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06922_ (.I(\mem.mem_dff.code_mem[10][5] ),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06923_ (.I(net238),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06924_ (.I(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06925_ (.A1(_02371_),
    .A2(_02367_),
    .B(_02361_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06926_ (.A1(_02369_),
    .A2(_02364_),
    .B(_02372_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06927_ (.I(\mem.mem_dff.code_mem[10][6] ),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06928_ (.A1(_02279_),
    .A2(_02367_),
    .B(_02361_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06929_ (.A1(_02373_),
    .A2(_02364_),
    .B(_02374_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06930_ (.I(\mem.mem_dff.code_mem[10][7] ),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06931_ (.I(_02127_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06932_ (.I(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06933_ (.I(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06934_ (.A1(_02282_),
    .A2(_02367_),
    .B(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06935_ (.A1(_02375_),
    .A2(_02364_),
    .B(_02379_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06936_ (.I(\mem.mem_dff.code_mem[11][0] ),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06937_ (.I(_02133_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06938_ (.A1(_02288_),
    .A2(_02319_),
    .A3(_02381_),
    .A4(_02135_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06939_ (.I(_02382_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_02286_),
    .A2(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06941_ (.I(_02384_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06942_ (.I(_02384_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06943_ (.A1(_02351_),
    .A2(_02386_),
    .B(_02378_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06944_ (.A1(_02380_),
    .A2(_02385_),
    .B(_02387_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06945_ (.I(\mem.mem_dff.code_mem[11][1] ),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06946_ (.I(_02143_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06947_ (.A1(_02389_),
    .A2(_02386_),
    .B(_02378_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06948_ (.A1(_02388_),
    .A2(_02385_),
    .B(_02390_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06949_ (.I(\mem.mem_dff.code_mem[11][2] ),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06950_ (.A1(_02358_),
    .A2(_02386_),
    .B(_02378_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06951_ (.A1(_02391_),
    .A2(_02385_),
    .B(_02392_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06952_ (.I(\mem.mem_dff.code_mem[11][3] ),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06953_ (.I(_02149_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06954_ (.I(_02377_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06955_ (.A1(_02394_),
    .A2(_02386_),
    .B(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06956_ (.A1(_02393_),
    .A2(_02385_),
    .B(_02396_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06957_ (.I(\mem.mem_dff.code_mem[11][4] ),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06958_ (.I(_02384_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06959_ (.I(_02384_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06960_ (.A1(_02366_),
    .A2(_02399_),
    .B(_02395_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06961_ (.A1(_02397_),
    .A2(_02398_),
    .B(_02400_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06962_ (.I(\mem.mem_dff.code_mem[11][5] ),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06963_ (.A1(_02371_),
    .A2(_02399_),
    .B(_02395_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06964_ (.A1(_02401_),
    .A2(_02398_),
    .B(_02402_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06965_ (.I(\mem.mem_dff.code_mem[11][6] ),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06966_ (.I(_02160_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06967_ (.A1(_02404_),
    .A2(_02399_),
    .B(_02395_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06968_ (.A1(_02403_),
    .A2(_02398_),
    .B(_02405_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06969_ (.I(\mem.mem_dff.code_mem[11][7] ),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06970_ (.I(_02164_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06971_ (.I(_02377_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06972_ (.A1(_02407_),
    .A2(_02399_),
    .B(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06973_ (.A1(_02406_),
    .A2(_02398_),
    .B(_02409_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06974_ (.I(\mem.mem_dff.code_mem[12][0] ),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06975_ (.I(_02017_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06976_ (.I(_02318_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06977_ (.A1(_02287_),
    .A2(_02412_),
    .A3(_02171_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06978_ (.I(_02413_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06979_ (.I(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(_02411_),
    .A2(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06981_ (.I(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06982_ (.I(_02416_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06983_ (.A1(_02351_),
    .A2(_02418_),
    .B(_02408_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06984_ (.A1(_02410_),
    .A2(_02417_),
    .B(_02419_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06985_ (.I(\mem.mem_dff.code_mem[12][1] ),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06986_ (.A1(_02389_),
    .A2(_02418_),
    .B(_02408_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06987_ (.A1(_02420_),
    .A2(_02417_),
    .B(_02421_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06988_ (.I(\mem.mem_dff.code_mem[12][2] ),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06989_ (.A1(_02358_),
    .A2(_02418_),
    .B(_02408_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06990_ (.A1(_02422_),
    .A2(_02417_),
    .B(_02423_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06991_ (.I(\mem.mem_dff.code_mem[12][3] ),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06992_ (.I(_02377_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06993_ (.A1(_02394_),
    .A2(_02418_),
    .B(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06994_ (.A1(_02424_),
    .A2(_02417_),
    .B(_02426_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06995_ (.I(\mem.mem_dff.code_mem[12][4] ),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06996_ (.I(_02416_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06997_ (.I(_02416_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06998_ (.A1(_02366_),
    .A2(_02429_),
    .B(_02425_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06999_ (.A1(_02427_),
    .A2(_02428_),
    .B(_02430_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07000_ (.I(\mem.mem_dff.code_mem[12][5] ),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07001_ (.A1(_02371_),
    .A2(_02429_),
    .B(_02425_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07002_ (.A1(_02431_),
    .A2(_02428_),
    .B(_02432_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07003_ (.I(\mem.mem_dff.code_mem[12][6] ),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07004_ (.A1(_02404_),
    .A2(_02429_),
    .B(_02425_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07005_ (.A1(_02433_),
    .A2(_02428_),
    .B(_02434_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07006_ (.I(\mem.mem_dff.code_mem[12][7] ),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07007_ (.I(_02376_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07008_ (.I(_02436_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07009_ (.A1(_02407_),
    .A2(_02429_),
    .B(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07010_ (.A1(_02435_),
    .A2(_02428_),
    .B(_02438_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07011_ (.I(\mem.mem_dff.code_mem[13][0] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07012_ (.I(_02318_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07013_ (.A1(_02345_),
    .A2(_02440_),
    .A3(_02198_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07014_ (.I(_02441_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07015_ (.I(_02442_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07016_ (.A1(_02411_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07017_ (.I(_02444_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07018_ (.I(_02444_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(_02351_),
    .A2(_02446_),
    .B(_02437_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07020_ (.A1(_02439_),
    .A2(_02445_),
    .B(_02447_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07021_ (.I(\mem.mem_dff.code_mem[13][1] ),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07022_ (.A1(_02389_),
    .A2(_02446_),
    .B(_02437_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07023_ (.A1(_02448_),
    .A2(_02445_),
    .B(_02449_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07024_ (.I(\mem.mem_dff.code_mem[13][2] ),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07025_ (.A1(_02358_),
    .A2(_02446_),
    .B(_02437_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07026_ (.A1(_02450_),
    .A2(_02445_),
    .B(_02451_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07027_ (.I(\mem.mem_dff.code_mem[13][3] ),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07028_ (.I(_02436_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07029_ (.A1(_02394_),
    .A2(_02446_),
    .B(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07030_ (.A1(_02452_),
    .A2(_02445_),
    .B(_02454_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07031_ (.I(\mem.mem_dff.code_mem[13][4] ),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07032_ (.I(_02444_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07033_ (.I(_02444_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07034_ (.A1(_02366_),
    .A2(_02457_),
    .B(_02453_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07035_ (.A1(_02455_),
    .A2(_02456_),
    .B(_02458_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07036_ (.I(\mem.mem_dff.code_mem[13][5] ),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07037_ (.A1(_02371_),
    .A2(_02457_),
    .B(_02453_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07038_ (.A1(_02459_),
    .A2(_02456_),
    .B(_02460_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07039_ (.I(\mem.mem_dff.code_mem[13][6] ),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07040_ (.A1(_02404_),
    .A2(_02457_),
    .B(_02453_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07041_ (.A1(_02461_),
    .A2(_02456_),
    .B(_02462_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07042_ (.I(\mem.mem_dff.code_mem[13][7] ),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07043_ (.I(_02436_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07044_ (.A1(_02407_),
    .A2(_02457_),
    .B(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07045_ (.A1(_02463_),
    .A2(_02456_),
    .B(_02465_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07046_ (.I(\mem.mem_dff.code_mem[14][0] ),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07047_ (.I(_02224_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07048_ (.A1(_02288_),
    .A2(_02319_),
    .A3(_02467_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07049_ (.I(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07050_ (.A1(_02411_),
    .A2(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07051_ (.I(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07052_ (.I(_02350_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07053_ (.I(_02470_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07054_ (.A1(_02472_),
    .A2(_02473_),
    .B(_02464_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07055_ (.A1(_02466_),
    .A2(_02471_),
    .B(_02474_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07056_ (.I(\mem.mem_dff.code_mem[14][1] ),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07057_ (.A1(_02389_),
    .A2(_02473_),
    .B(_02464_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07058_ (.A1(_02475_),
    .A2(_02471_),
    .B(_02476_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07059_ (.I(\mem.mem_dff.code_mem[14][2] ),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07060_ (.I(_02357_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07061_ (.A1(_02478_),
    .A2(_02473_),
    .B(_02464_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07062_ (.A1(_02477_),
    .A2(_02471_),
    .B(_02479_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07063_ (.I(\mem.mem_dff.code_mem[14][3] ),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07064_ (.I(_02436_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07065_ (.A1(_02394_),
    .A2(_02473_),
    .B(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07066_ (.A1(_02480_),
    .A2(_02471_),
    .B(_02482_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07067_ (.I(\mem.mem_dff.code_mem[14][4] ),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07068_ (.I(_02470_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07069_ (.I(_02365_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07070_ (.I(_02470_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07071_ (.A1(_02485_),
    .A2(_02486_),
    .B(_02481_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07072_ (.A1(_02483_),
    .A2(_02484_),
    .B(_02487_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07073_ (.I(\mem.mem_dff.code_mem[14][5] ),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07074_ (.I(_02370_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07075_ (.A1(_02489_),
    .A2(_02486_),
    .B(_02481_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07076_ (.A1(_02488_),
    .A2(_02484_),
    .B(_02490_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07077_ (.I(\mem.mem_dff.code_mem[14][6] ),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07078_ (.A1(_02404_),
    .A2(_02486_),
    .B(_02481_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07079_ (.A1(_02491_),
    .A2(_02484_),
    .B(_02492_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07080_ (.I(\mem.mem_dff.code_mem[14][7] ),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07081_ (.I(_02376_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07082_ (.I(_02494_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07083_ (.A1(_02407_),
    .A2(_02486_),
    .B(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07084_ (.A1(_02493_),
    .A2(_02484_),
    .B(_02496_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07085_ (.I(\mem.mem_dff.code_mem[15][0] ),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07086_ (.A1(_02287_),
    .A2(_02412_),
    .A3(_02255_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07087_ (.I(_02498_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07088_ (.A1(_02411_),
    .A2(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07089_ (.I(_02500_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07090_ (.I(_02500_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07091_ (.A1(_02472_),
    .A2(_02502_),
    .B(_02495_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07092_ (.A1(_02497_),
    .A2(_02501_),
    .B(_02503_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07093_ (.I(\mem.mem_dff.code_mem[15][1] ),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07094_ (.I(_02036_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07095_ (.I(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07096_ (.A1(_02506_),
    .A2(_02502_),
    .B(_02495_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07097_ (.A1(_02504_),
    .A2(_02501_),
    .B(_02507_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07098_ (.I(\mem.mem_dff.code_mem[15][2] ),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07099_ (.A1(_02478_),
    .A2(_02502_),
    .B(_02495_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07100_ (.A1(_02508_),
    .A2(_02501_),
    .B(_02509_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07101_ (.I(\mem.mem_dff.code_mem[15][3] ),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07102_ (.I(_02044_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07103_ (.I(_02511_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07104_ (.I(_02494_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07105_ (.A1(_02512_),
    .A2(_02502_),
    .B(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07106_ (.A1(_02510_),
    .A2(_02501_),
    .B(_02514_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07107_ (.I(\mem.mem_dff.code_mem[15][4] ),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07108_ (.I(_02500_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07109_ (.I(_02500_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07110_ (.A1(_02485_),
    .A2(_02517_),
    .B(_02513_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07111_ (.A1(_02515_),
    .A2(_02516_),
    .B(_02518_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07112_ (.I(\mem.mem_dff.code_mem[15][5] ),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07113_ (.A1(_02489_),
    .A2(_02517_),
    .B(_02513_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07114_ (.A1(_02519_),
    .A2(_02516_),
    .B(_02520_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07115_ (.I(\mem.mem_dff.code_mem[15][6] ),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07116_ (.I(_02059_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07117_ (.I(_02522_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07118_ (.A1(_02523_),
    .A2(_02517_),
    .B(_02513_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07119_ (.A1(_02521_),
    .A2(_02516_),
    .B(_02524_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07120_ (.I(\mem.mem_dff.code_mem[15][7] ),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07121_ (.I(_02063_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07122_ (.I(_02526_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07123_ (.I(_02494_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07124_ (.A1(_02527_),
    .A2(_02517_),
    .B(_02528_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07125_ (.A1(_02525_),
    .A2(_02516_),
    .B(_02529_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07126_ (.I(\mem.mem_dff.code_mem[16][0] ),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07127_ (.I(_02016_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07128_ (.I(_02531_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07129_ (.A1(net187),
    .A2(_02023_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07130_ (.I(_02533_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07131_ (.A1(_02021_),
    .A2(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07132_ (.I(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07133_ (.A1(_02532_),
    .A2(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07134_ (.I(_02537_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07135_ (.I(_02537_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07136_ (.A1(_02472_),
    .A2(_02539_),
    .B(_02528_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07137_ (.A1(_02530_),
    .A2(_02538_),
    .B(_02540_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07138_ (.I(\mem.mem_dff.code_mem[16][1] ),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07139_ (.A1(_02506_),
    .A2(_02539_),
    .B(_02528_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07140_ (.A1(_02541_),
    .A2(_02538_),
    .B(_02542_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07141_ (.I(\mem.mem_dff.code_mem[16][2] ),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07142_ (.A1(_02478_),
    .A2(_02539_),
    .B(_02528_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07143_ (.A1(_02543_),
    .A2(_02538_),
    .B(_02544_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07144_ (.I(\mem.mem_dff.code_mem[16][3] ),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07145_ (.I(_02494_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07146_ (.A1(_02512_),
    .A2(_02539_),
    .B(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07147_ (.A1(_02545_),
    .A2(_02538_),
    .B(_02547_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07148_ (.I(\mem.mem_dff.code_mem[16][4] ),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07149_ (.I(_02537_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07150_ (.I(_02537_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07151_ (.A1(_02485_),
    .A2(_02550_),
    .B(_02546_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07152_ (.A1(_02548_),
    .A2(_02549_),
    .B(_02551_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07153_ (.I(\mem.mem_dff.code_mem[16][5] ),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07154_ (.A1(_02489_),
    .A2(_02550_),
    .B(_02546_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07155_ (.A1(_02552_),
    .A2(_02549_),
    .B(_02553_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07156_ (.I(\mem.mem_dff.code_mem[16][6] ),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07157_ (.A1(_02523_),
    .A2(_02550_),
    .B(_02546_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07158_ (.A1(_02554_),
    .A2(_02549_),
    .B(_02555_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07159_ (.I(\mem.mem_dff.code_mem[16][7] ),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07160_ (.I(_02376_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07161_ (.I(_02557_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07162_ (.A1(_02527_),
    .A2(_02550_),
    .B(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07163_ (.A1(_02556_),
    .A2(_02549_),
    .B(_02559_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07164_ (.I(\mem.mem_dff.code_mem[17][0] ),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07165_ (.A1(_02069_),
    .A2(_02534_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07166_ (.I(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07167_ (.A1(_02532_),
    .A2(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07168_ (.I(_02563_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07169_ (.I(_02563_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07170_ (.A1(_02472_),
    .A2(_02565_),
    .B(_02558_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07171_ (.A1(_02560_),
    .A2(_02564_),
    .B(_02566_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07172_ (.I(\mem.mem_dff.code_mem[17][1] ),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07173_ (.A1(_02506_),
    .A2(_02565_),
    .B(_02558_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07174_ (.A1(_02567_),
    .A2(_02564_),
    .B(_02568_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07175_ (.I(\mem.mem_dff.code_mem[17][2] ),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07176_ (.A1(_02478_),
    .A2(_02565_),
    .B(_02558_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07177_ (.A1(_02569_),
    .A2(_02564_),
    .B(_02570_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07178_ (.I(\mem.mem_dff.code_mem[17][3] ),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07179_ (.I(_02557_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07180_ (.A1(_02512_),
    .A2(_02565_),
    .B(_02572_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07181_ (.A1(_02571_),
    .A2(_02564_),
    .B(_02573_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07182_ (.I(\mem.mem_dff.code_mem[17][4] ),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07183_ (.I(_02563_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07184_ (.I(_02563_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07185_ (.A1(_02485_),
    .A2(_02576_),
    .B(_02572_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07186_ (.A1(_02574_),
    .A2(_02575_),
    .B(_02577_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07187_ (.I(\mem.mem_dff.code_mem[17][5] ),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07188_ (.A1(_02489_),
    .A2(_02576_),
    .B(_02572_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07189_ (.A1(_02578_),
    .A2(_02575_),
    .B(_02579_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07190_ (.I(\mem.mem_dff.code_mem[17][6] ),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07191_ (.A1(_02523_),
    .A2(_02576_),
    .B(_02572_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07192_ (.A1(_02580_),
    .A2(_02575_),
    .B(_02581_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07193_ (.I(\mem.mem_dff.code_mem[17][7] ),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07194_ (.I(_02557_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07195_ (.A1(_02527_),
    .A2(_02576_),
    .B(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07196_ (.A1(_02582_),
    .A2(_02575_),
    .B(_02584_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07197_ (.I(\mem.mem_dff.code_mem[18][0] ),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07198_ (.I(_02533_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07199_ (.A1(_02096_),
    .A2(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07200_ (.I(_02587_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(_02532_),
    .A2(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07202_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07203_ (.I(_02350_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07204_ (.I(_02589_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07205_ (.A1(_02591_),
    .A2(_02592_),
    .B(_02583_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07206_ (.A1(_02585_),
    .A2(_02590_),
    .B(_02593_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07207_ (.I(\mem.mem_dff.code_mem[18][1] ),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07208_ (.A1(_02506_),
    .A2(_02592_),
    .B(_02583_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07209_ (.A1(_02594_),
    .A2(_02590_),
    .B(_02595_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07210_ (.I(\mem.mem_dff.code_mem[18][2] ),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07211_ (.I(_02357_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07212_ (.A1(_02597_),
    .A2(_02592_),
    .B(_02583_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07213_ (.A1(_02596_),
    .A2(_02590_),
    .B(_02598_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07214_ (.I(\mem.mem_dff.code_mem[18][3] ),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07215_ (.I(_02557_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07216_ (.A1(_02512_),
    .A2(_02592_),
    .B(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07217_ (.A1(_02599_),
    .A2(_02590_),
    .B(_02601_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07218_ (.I(\mem.mem_dff.code_mem[18][4] ),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07219_ (.I(_02589_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07220_ (.I(_02365_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07221_ (.I(_02589_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(_02604_),
    .A2(_02605_),
    .B(_02600_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07223_ (.A1(_02602_),
    .A2(_02603_),
    .B(_02606_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07224_ (.I(\mem.mem_dff.code_mem[18][5] ),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07225_ (.I(_02370_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07226_ (.A1(_02608_),
    .A2(_02605_),
    .B(_02600_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07227_ (.A1(_02607_),
    .A2(_02603_),
    .B(_02609_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07228_ (.I(\mem.mem_dff.code_mem[18][6] ),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07229_ (.A1(_02523_),
    .A2(_02605_),
    .B(_02600_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07230_ (.A1(_02610_),
    .A2(_02603_),
    .B(_02611_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07231_ (.I(\mem.mem_dff.code_mem[18][7] ),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07232_ (.I(_02127_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07233_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07234_ (.I(_02614_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07235_ (.A1(_02527_),
    .A2(_02605_),
    .B(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07236_ (.A1(_02612_),
    .A2(_02603_),
    .B(_02616_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07237_ (.I(\mem.mem_dff.code_mem[19][0] ),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07238_ (.I(_00760_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07239_ (.A1(_02133_),
    .A2(_02618_),
    .A3(_02586_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07240_ (.I(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07241_ (.A1(_02532_),
    .A2(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07242_ (.I(_02621_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07243_ (.I(_02621_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07244_ (.A1(_02591_),
    .A2(_02623_),
    .B(_02615_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07245_ (.A1(_02617_),
    .A2(_02622_),
    .B(_02624_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07246_ (.I(\mem.mem_dff.code_mem[19][1] ),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07247_ (.I(_02505_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07248_ (.A1(_02626_),
    .A2(_02623_),
    .B(_02615_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07249_ (.A1(_02625_),
    .A2(_02622_),
    .B(_02627_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07250_ (.I(\mem.mem_dff.code_mem[19][2] ),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07251_ (.A1(_02597_),
    .A2(_02623_),
    .B(_02615_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07252_ (.A1(_02628_),
    .A2(_02622_),
    .B(_02629_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07253_ (.I(\mem.mem_dff.code_mem[19][3] ),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07254_ (.I(_02511_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07255_ (.I(_02614_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07256_ (.A1(_02631_),
    .A2(_02623_),
    .B(_02632_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07257_ (.A1(_02630_),
    .A2(_02622_),
    .B(_02633_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07258_ (.I(\mem.mem_dff.code_mem[19][4] ),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07259_ (.I(_02621_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07260_ (.I(_02621_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07261_ (.A1(_02604_),
    .A2(_02636_),
    .B(_02632_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07262_ (.A1(_02634_),
    .A2(_02635_),
    .B(_02637_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07263_ (.I(\mem.mem_dff.code_mem[19][5] ),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07264_ (.A1(_02608_),
    .A2(_02636_),
    .B(_02632_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07265_ (.A1(_02638_),
    .A2(_02635_),
    .B(_02639_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07266_ (.I(\mem.mem_dff.code_mem[19][6] ),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07267_ (.I(_02522_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07268_ (.A1(_02641_),
    .A2(_02636_),
    .B(_02632_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07269_ (.A1(_02640_),
    .A2(_02635_),
    .B(_02642_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07270_ (.I(\mem.mem_dff.code_mem[19][7] ),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07271_ (.I(_02526_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07272_ (.I(_02614_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07273_ (.A1(_02644_),
    .A2(_02636_),
    .B(_02645_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07274_ (.A1(_02643_),
    .A2(_02635_),
    .B(_02646_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07275_ (.I(\mem.mem_dff.code_mem[20][0] ),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07276_ (.I(_02531_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07277_ (.A1(_02171_),
    .A2(_02534_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07278_ (.I(_02649_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07279_ (.A1(_02648_),
    .A2(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07280_ (.I(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07281_ (.I(_02651_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07282_ (.A1(_02591_),
    .A2(_02653_),
    .B(_02645_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07283_ (.A1(_02647_),
    .A2(_02652_),
    .B(_02654_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07284_ (.I(\mem.mem_dff.code_mem[20][1] ),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07285_ (.A1(_02626_),
    .A2(_02653_),
    .B(_02645_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07286_ (.A1(_02655_),
    .A2(_02652_),
    .B(_02656_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07287_ (.I(\mem.mem_dff.code_mem[20][2] ),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07288_ (.A1(_02597_),
    .A2(_02653_),
    .B(_02645_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07289_ (.A1(_02657_),
    .A2(_02652_),
    .B(_02658_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07290_ (.I(\mem.mem_dff.code_mem[20][3] ),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07291_ (.I(_02614_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07292_ (.A1(_02631_),
    .A2(_02653_),
    .B(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07293_ (.A1(_02659_),
    .A2(_02652_),
    .B(_02661_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07294_ (.I(\mem.mem_dff.code_mem[20][4] ),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07295_ (.I(_02651_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07296_ (.I(_02651_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07297_ (.A1(_02604_),
    .A2(_02664_),
    .B(_02660_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07298_ (.A1(_02662_),
    .A2(_02663_),
    .B(_02665_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07299_ (.I(\mem.mem_dff.code_mem[20][5] ),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07300_ (.A1(_02608_),
    .A2(_02664_),
    .B(_02660_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07301_ (.A1(_02666_),
    .A2(_02663_),
    .B(_02667_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07302_ (.I(\mem.mem_dff.code_mem[20][6] ),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07303_ (.A1(_02641_),
    .A2(_02664_),
    .B(_02660_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07304_ (.A1(_02668_),
    .A2(_02663_),
    .B(_02669_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07305_ (.I(\mem.mem_dff.code_mem[20][7] ),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07306_ (.I(_02613_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07307_ (.I(_02671_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07308_ (.A1(_02644_),
    .A2(_02664_),
    .B(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07309_ (.A1(_02670_),
    .A2(_02663_),
    .B(_02673_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07310_ (.I(\mem.mem_dff.code_mem[21][0] ),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07311_ (.A1(_02198_),
    .A2(_02586_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07312_ (.I(_02675_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07313_ (.A1(_02648_),
    .A2(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07314_ (.I(_02677_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07315_ (.I(_02677_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07316_ (.A1(_02591_),
    .A2(_02679_),
    .B(_02672_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07317_ (.A1(_02674_),
    .A2(_02678_),
    .B(_02680_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07318_ (.I(\mem.mem_dff.code_mem[21][1] ),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07319_ (.A1(_02626_),
    .A2(_02679_),
    .B(_02672_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07320_ (.A1(_02681_),
    .A2(_02678_),
    .B(_02682_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07321_ (.I(\mem.mem_dff.code_mem[21][2] ),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07322_ (.A1(_02597_),
    .A2(_02679_),
    .B(_02672_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07323_ (.A1(_02683_),
    .A2(_02678_),
    .B(_02684_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07324_ (.I(\mem.mem_dff.code_mem[21][3] ),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07325_ (.I(_02671_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07326_ (.A1(_02631_),
    .A2(_02679_),
    .B(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07327_ (.A1(_02685_),
    .A2(_02678_),
    .B(_02687_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07328_ (.I(\mem.mem_dff.code_mem[21][4] ),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07329_ (.I(_02677_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07330_ (.I(_02677_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07331_ (.A1(_02604_),
    .A2(_02690_),
    .B(_02686_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07332_ (.A1(_02688_),
    .A2(_02689_),
    .B(_02691_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07333_ (.I(\mem.mem_dff.code_mem[21][5] ),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07334_ (.A1(_02608_),
    .A2(_02690_),
    .B(_02686_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07335_ (.A1(_02692_),
    .A2(_02689_),
    .B(_02693_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07336_ (.I(\mem.mem_dff.code_mem[21][6] ),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07337_ (.A1(_02641_),
    .A2(_02690_),
    .B(_02686_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07338_ (.A1(_02694_),
    .A2(_02689_),
    .B(_02695_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07339_ (.I(\mem.mem_dff.code_mem[21][7] ),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07340_ (.I(_02671_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07341_ (.A1(_02644_),
    .A2(_02690_),
    .B(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07342_ (.A1(_02696_),
    .A2(_02689_),
    .B(_02698_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07343_ (.I(\mem.mem_dff.code_mem[22][0] ),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07344_ (.A1(_02467_),
    .A2(_02534_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07345_ (.I(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07346_ (.A1(_02648_),
    .A2(_02701_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07347_ (.I(_02702_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07348_ (.I(_02350_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07349_ (.I(_02702_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07350_ (.A1(_02704_),
    .A2(_02705_),
    .B(_02697_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07351_ (.A1(_02699_),
    .A2(_02703_),
    .B(_02706_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07352_ (.I(\mem.mem_dff.code_mem[22][1] ),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07353_ (.A1(_02626_),
    .A2(_02705_),
    .B(_02697_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07354_ (.A1(_02707_),
    .A2(_02703_),
    .B(_02708_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07355_ (.I(\mem.mem_dff.code_mem[22][2] ),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07356_ (.I(_02357_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(_02710_),
    .A2(_02705_),
    .B(_02697_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07358_ (.A1(_02709_),
    .A2(_02703_),
    .B(_02711_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07359_ (.I(\mem.mem_dff.code_mem[22][3] ),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07360_ (.I(_02671_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07361_ (.A1(_02631_),
    .A2(_02705_),
    .B(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07362_ (.A1(_02712_),
    .A2(_02703_),
    .B(_02714_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07363_ (.I(\mem.mem_dff.code_mem[22][4] ),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07364_ (.I(_02702_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07365_ (.I(_02365_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07366_ (.I(_02702_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(_02717_),
    .A2(_02718_),
    .B(_02713_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07368_ (.A1(_02715_),
    .A2(_02716_),
    .B(_02719_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07369_ (.I(\mem.mem_dff.code_mem[22][5] ),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07370_ (.I(_02370_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07371_ (.A1(_02721_),
    .A2(_02718_),
    .B(_02713_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07372_ (.A1(_02720_),
    .A2(_02716_),
    .B(_02722_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07373_ (.I(\mem.mem_dff.code_mem[22][6] ),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07374_ (.A1(_02641_),
    .A2(_02718_),
    .B(_02713_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07375_ (.A1(_02723_),
    .A2(_02716_),
    .B(_02724_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07376_ (.I(\mem.mem_dff.code_mem[22][7] ),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07377_ (.I(_02613_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07378_ (.I(_02726_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07379_ (.A1(_02644_),
    .A2(_02718_),
    .B(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07380_ (.A1(_02725_),
    .A2(_02716_),
    .B(_02728_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07381_ (.I(\mem.mem_dff.code_mem[23][0] ),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07382_ (.A1(_02255_),
    .A2(_02586_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07383_ (.I(_02730_),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07384_ (.A1(_02648_),
    .A2(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07385_ (.I(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07386_ (.I(_02732_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07387_ (.A1(_02704_),
    .A2(_02734_),
    .B(_02727_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07388_ (.A1(_02729_),
    .A2(_02733_),
    .B(_02735_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07389_ (.I(\mem.mem_dff.code_mem[23][1] ),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07390_ (.I(_02505_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07391_ (.A1(_02737_),
    .A2(_02734_),
    .B(_02727_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07392_ (.A1(_02736_),
    .A2(_02733_),
    .B(_02738_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07393_ (.I(\mem.mem_dff.code_mem[23][2] ),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07394_ (.A1(_02710_),
    .A2(_02734_),
    .B(_02727_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07395_ (.A1(_02739_),
    .A2(_02733_),
    .B(_02740_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07396_ (.I(\mem.mem_dff.code_mem[23][3] ),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07397_ (.I(_02511_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07398_ (.I(_02726_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07399_ (.A1(_02742_),
    .A2(_02734_),
    .B(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07400_ (.A1(_02741_),
    .A2(_02733_),
    .B(_02744_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07401_ (.I(\mem.mem_dff.code_mem[23][4] ),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07402_ (.I(_02732_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07403_ (.I(_02732_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07404_ (.A1(_02717_),
    .A2(_02747_),
    .B(_02743_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07405_ (.A1(_02745_),
    .A2(_02746_),
    .B(_02748_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07406_ (.I(\mem.mem_dff.code_mem[23][5] ),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07407_ (.A1(_02721_),
    .A2(_02747_),
    .B(_02743_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07408_ (.A1(_02749_),
    .A2(_02746_),
    .B(_02750_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07409_ (.I(\mem.mem_dff.code_mem[23][6] ),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07410_ (.I(_02522_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07411_ (.A1(_02752_),
    .A2(_02747_),
    .B(_02743_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07412_ (.A1(_02751_),
    .A2(_02746_),
    .B(_02753_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07413_ (.I(\mem.mem_dff.code_mem[23][7] ),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07414_ (.I(_02526_),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07415_ (.I(_02726_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07416_ (.A1(_02755_),
    .A2(_02747_),
    .B(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07417_ (.A1(_02754_),
    .A2(_02746_),
    .B(_02757_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07418_ (.I(\mem.mem_dff.code_mem[24][0] ),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07419_ (.I(_02531_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07420_ (.I(_02022_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07421_ (.A1(_02760_),
    .A2(_02291_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07422_ (.I(_02761_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(_02759_),
    .A2(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07424_ (.I(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07425_ (.I(_02763_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07426_ (.A1(_02704_),
    .A2(_02765_),
    .B(_02756_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07427_ (.A1(_02758_),
    .A2(_02764_),
    .B(_02766_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07428_ (.I(\mem.mem_dff.code_mem[24][1] ),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07429_ (.A1(_02737_),
    .A2(_02765_),
    .B(_02756_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07430_ (.A1(_02767_),
    .A2(_02764_),
    .B(_02768_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07431_ (.I(\mem.mem_dff.code_mem[24][2] ),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07432_ (.A1(_02710_),
    .A2(_02765_),
    .B(_02756_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07433_ (.A1(_02769_),
    .A2(_02764_),
    .B(_02770_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07434_ (.I(\mem.mem_dff.code_mem[24][3] ),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07435_ (.I(_02726_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07436_ (.A1(_02742_),
    .A2(_02765_),
    .B(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07437_ (.A1(_02771_),
    .A2(_02764_),
    .B(_02773_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07438_ (.I(\mem.mem_dff.code_mem[24][4] ),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07439_ (.I(_02763_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07440_ (.I(_02763_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07441_ (.A1(_02717_),
    .A2(_02776_),
    .B(_02772_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07442_ (.A1(_02774_),
    .A2(_02775_),
    .B(_02777_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07443_ (.I(\mem.mem_dff.code_mem[24][5] ),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07444_ (.A1(_02721_),
    .A2(_02776_),
    .B(_02772_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07445_ (.A1(_02778_),
    .A2(_02775_),
    .B(_02779_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07446_ (.I(\mem.mem_dff.code_mem[24][6] ),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07447_ (.A1(_02752_),
    .A2(_02776_),
    .B(_02772_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07448_ (.A1(_02780_),
    .A2(_02775_),
    .B(_02781_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07449_ (.I(\mem.mem_dff.code_mem[24][7] ),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07450_ (.I(_02613_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07451_ (.I(_02783_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07452_ (.A1(_02755_),
    .A2(_02776_),
    .B(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07453_ (.A1(_02782_),
    .A2(_02775_),
    .B(_02785_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07454_ (.I(\mem.mem_dff.code_mem[25][0] ),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07455_ (.I(_02022_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07456_ (.A1(_02787_),
    .A2(_02440_),
    .A3(_02069_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07457_ (.I(_02788_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(_02759_),
    .A2(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07459_ (.I(_02790_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07460_ (.I(_02790_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07461_ (.A1(_02704_),
    .A2(_02792_),
    .B(_02784_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07462_ (.A1(_02786_),
    .A2(_02791_),
    .B(_02793_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07463_ (.I(\mem.mem_dff.code_mem[25][1] ),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07464_ (.A1(_02737_),
    .A2(_02792_),
    .B(_02784_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07465_ (.A1(_02794_),
    .A2(_02791_),
    .B(_02795_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07466_ (.I(\mem.mem_dff.code_mem[25][2] ),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07467_ (.A1(_02710_),
    .A2(_02792_),
    .B(_02784_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07468_ (.A1(_02796_),
    .A2(_02791_),
    .B(_02797_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07469_ (.I(\mem.mem_dff.code_mem[25][3] ),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07470_ (.I(_02783_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07471_ (.A1(_02742_),
    .A2(_02792_),
    .B(_02799_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07472_ (.A1(_02798_),
    .A2(_02791_),
    .B(_02800_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07473_ (.I(\mem.mem_dff.code_mem[25][4] ),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07474_ (.I(_02790_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07475_ (.I(_02790_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07476_ (.A1(_02717_),
    .A2(_02803_),
    .B(_02799_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07477_ (.A1(_02801_),
    .A2(_02802_),
    .B(_02804_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07478_ (.I(\mem.mem_dff.code_mem[25][5] ),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07479_ (.A1(_02721_),
    .A2(_02803_),
    .B(_02799_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07480_ (.A1(_02805_),
    .A2(_02802_),
    .B(_02806_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07481_ (.I(\mem.mem_dff.code_mem[25][6] ),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07482_ (.A1(_02752_),
    .A2(_02803_),
    .B(_02799_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07483_ (.A1(_02807_),
    .A2(_02802_),
    .B(_02808_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07484_ (.I(\mem.mem_dff.code_mem[25][7] ),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07485_ (.I(_02783_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07486_ (.A1(_02755_),
    .A2(_02803_),
    .B(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07487_ (.A1(_02809_),
    .A2(_02802_),
    .B(_02811_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07488_ (.I(\mem.mem_dff.code_mem[26][0] ),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07489_ (.I(_02412_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07490_ (.A1(_02760_),
    .A2(_02813_),
    .A3(_02096_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07491_ (.I(_02814_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07492_ (.A1(_02759_),
    .A2(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07493_ (.I(_02816_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07494_ (.I(_02030_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07495_ (.I(_02816_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07496_ (.A1(_02818_),
    .A2(_02819_),
    .B(_02810_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07497_ (.A1(_02812_),
    .A2(_02817_),
    .B(_02820_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07498_ (.I(\mem.mem_dff.code_mem[26][1] ),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07499_ (.A1(_02737_),
    .A2(_02819_),
    .B(_02810_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07500_ (.A1(_02821_),
    .A2(_02817_),
    .B(_02822_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07501_ (.I(\mem.mem_dff.code_mem[26][2] ),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07502_ (.I(_02040_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07503_ (.A1(_02824_),
    .A2(_02819_),
    .B(_02810_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07504_ (.A1(_02823_),
    .A2(_02817_),
    .B(_02825_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07505_ (.I(\mem.mem_dff.code_mem[26][3] ),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07506_ (.I(_02783_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07507_ (.A1(_02742_),
    .A2(_02819_),
    .B(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07508_ (.A1(_02826_),
    .A2(_02817_),
    .B(_02828_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07509_ (.I(\mem.mem_dff.code_mem[26][4] ),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07510_ (.I(_02816_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07511_ (.I(_02050_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07512_ (.I(_02816_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07513_ (.A1(_02831_),
    .A2(_02832_),
    .B(_02827_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07514_ (.A1(_02829_),
    .A2(_02830_),
    .B(_02833_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07515_ (.I(\mem.mem_dff.code_mem[26][5] ),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07516_ (.I(_02055_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07517_ (.A1(_02835_),
    .A2(_02832_),
    .B(_02827_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07518_ (.A1(_02834_),
    .A2(_02830_),
    .B(_02836_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07519_ (.I(\mem.mem_dff.code_mem[26][6] ),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07520_ (.A1(_02752_),
    .A2(_02832_),
    .B(_02827_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07521_ (.A1(_02837_),
    .A2(_02830_),
    .B(_02838_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07522_ (.I(\mem.mem_dff.code_mem[26][7] ),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07523_ (.I(_01997_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07524_ (.I(_02840_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07525_ (.I(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07526_ (.A1(_02755_),
    .A2(_02832_),
    .B(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07527_ (.A1(_02839_),
    .A2(_02830_),
    .B(_02843_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07528_ (.I(\mem.mem_dff.code_mem[27][0] ),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07529_ (.A1(_02022_),
    .A2(_02318_),
    .A3(_02133_),
    .A4(_02618_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07530_ (.I(_02845_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(_02759_),
    .A2(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07532_ (.I(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07533_ (.I(_02847_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07534_ (.A1(_02818_),
    .A2(_02849_),
    .B(_02842_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07535_ (.A1(_02844_),
    .A2(_02848_),
    .B(_02850_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07536_ (.I(\mem.mem_dff.code_mem[27][1] ),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07537_ (.I(_02505_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07538_ (.A1(_02852_),
    .A2(_02849_),
    .B(_02842_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07539_ (.A1(_02851_),
    .A2(_02848_),
    .B(_02853_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07540_ (.I(\mem.mem_dff.code_mem[27][2] ),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07541_ (.A1(_02824_),
    .A2(_02849_),
    .B(_02842_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07542_ (.A1(_02854_),
    .A2(_02848_),
    .B(_02855_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07543_ (.I(\mem.mem_dff.code_mem[27][3] ),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07544_ (.I(_02511_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07545_ (.I(_02841_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07546_ (.A1(_02857_),
    .A2(_02849_),
    .B(_02858_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07547_ (.A1(_02856_),
    .A2(_02848_),
    .B(_02859_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07548_ (.I(\mem.mem_dff.code_mem[27][4] ),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07549_ (.I(_02847_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07550_ (.I(_02847_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07551_ (.A1(_02831_),
    .A2(_02862_),
    .B(_02858_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07552_ (.A1(_02860_),
    .A2(_02861_),
    .B(_02863_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07553_ (.I(\mem.mem_dff.code_mem[27][5] ),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07554_ (.A1(_02835_),
    .A2(_02862_),
    .B(_02858_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07555_ (.A1(_02864_),
    .A2(_02861_),
    .B(_02865_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07556_ (.I(\mem.mem_dff.code_mem[27][6] ),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07557_ (.I(_02522_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07558_ (.A1(_02867_),
    .A2(_02862_),
    .B(_02858_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07559_ (.A1(_02866_),
    .A2(_02861_),
    .B(_02868_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07560_ (.I(\mem.mem_dff.code_mem[27][7] ),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07561_ (.I(_02526_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07562_ (.I(_02841_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07563_ (.A1(_02870_),
    .A2(_02862_),
    .B(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07564_ (.A1(_02869_),
    .A2(_02861_),
    .B(_02872_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07565_ (.I(\mem.mem_dff.code_mem[28][0] ),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07566_ (.I(_02531_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07567_ (.A1(_02760_),
    .A2(_02813_),
    .A3(_02171_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07568_ (.I(_02875_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(_02874_),
    .A2(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07570_ (.I(_02877_),
    .Z(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07571_ (.I(_02877_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07572_ (.A1(_02818_),
    .A2(_02879_),
    .B(_02871_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07573_ (.A1(_02873_),
    .A2(_02878_),
    .B(_02880_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07574_ (.I(\mem.mem_dff.code_mem[28][1] ),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07575_ (.A1(_02852_),
    .A2(_02879_),
    .B(_02871_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07576_ (.A1(_02881_),
    .A2(_02878_),
    .B(_02882_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07577_ (.I(\mem.mem_dff.code_mem[28][2] ),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07578_ (.A1(_02824_),
    .A2(_02879_),
    .B(_02871_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07579_ (.A1(_02883_),
    .A2(_02878_),
    .B(_02884_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07580_ (.I(\mem.mem_dff.code_mem[28][3] ),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07581_ (.I(_02841_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07582_ (.A1(_02857_),
    .A2(_02879_),
    .B(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07583_ (.A1(_02885_),
    .A2(_02878_),
    .B(_02887_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07584_ (.I(\mem.mem_dff.code_mem[28][4] ),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07585_ (.I(_02877_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07586_ (.I(_02877_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07587_ (.A1(_02831_),
    .A2(_02890_),
    .B(_02886_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07588_ (.A1(_02888_),
    .A2(_02889_),
    .B(_02891_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07589_ (.I(\mem.mem_dff.code_mem[28][5] ),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07590_ (.A1(_02835_),
    .A2(_02890_),
    .B(_02886_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07591_ (.A1(_02892_),
    .A2(_02889_),
    .B(_02893_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07592_ (.I(\mem.mem_dff.code_mem[28][6] ),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07593_ (.A1(_02867_),
    .A2(_02890_),
    .B(_02886_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07594_ (.A1(_02894_),
    .A2(_02889_),
    .B(_02895_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07595_ (.I(\mem.mem_dff.code_mem[28][7] ),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07596_ (.I(_02840_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07597_ (.I(_02897_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07598_ (.A1(_02870_),
    .A2(_02890_),
    .B(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07599_ (.A1(_02896_),
    .A2(_02889_),
    .B(_02899_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07600_ (.I(\mem.mem_dff.code_mem[29][0] ),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07601_ (.A1(_02787_),
    .A2(_02440_),
    .A3(_02198_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07602_ (.I(_02901_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07603_ (.A1(_02874_),
    .A2(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07604_ (.I(_02903_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07605_ (.I(_02903_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07606_ (.A1(_02818_),
    .A2(_02905_),
    .B(_02898_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07607_ (.A1(_02900_),
    .A2(_02904_),
    .B(_02906_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07608_ (.I(\mem.mem_dff.code_mem[29][1] ),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07609_ (.A1(_02852_),
    .A2(_02905_),
    .B(_02898_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07610_ (.A1(_02907_),
    .A2(_02904_),
    .B(_02908_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07611_ (.I(\mem.mem_dff.code_mem[29][2] ),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07612_ (.A1(_02824_),
    .A2(_02905_),
    .B(_02898_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07613_ (.A1(_02909_),
    .A2(_02904_),
    .B(_02910_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07614_ (.I(\mem.mem_dff.code_mem[29][3] ),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07615_ (.I(_02897_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07616_ (.A1(_02857_),
    .A2(_02905_),
    .B(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07617_ (.A1(_02911_),
    .A2(_02904_),
    .B(_02913_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07618_ (.I(\mem.mem_dff.code_mem[29][4] ),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07619_ (.I(_02903_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07620_ (.I(_02903_),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07621_ (.A1(_02831_),
    .A2(_02916_),
    .B(_02912_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07622_ (.A1(_02914_),
    .A2(_02915_),
    .B(_02917_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07623_ (.I(\mem.mem_dff.code_mem[29][5] ),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07624_ (.A1(_02835_),
    .A2(_02916_),
    .B(_02912_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07625_ (.A1(_02918_),
    .A2(_02915_),
    .B(_02919_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07626_ (.I(\mem.mem_dff.code_mem[29][6] ),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07627_ (.A1(_02867_),
    .A2(_02916_),
    .B(_02912_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07628_ (.A1(_02920_),
    .A2(_02915_),
    .B(_02921_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07629_ (.I(\mem.mem_dff.code_mem[29][7] ),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07630_ (.I(_02897_),
    .Z(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07631_ (.A1(_02870_),
    .A2(_02916_),
    .B(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07632_ (.A1(_02922_),
    .A2(_02915_),
    .B(_02924_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07633_ (.I(\mem.mem_dff.code_mem[30][0] ),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07634_ (.A1(_02787_),
    .A2(_02440_),
    .A3(_02224_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07635_ (.I(_02926_),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07636_ (.A1(_02874_),
    .A2(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07637_ (.I(_02928_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07638_ (.I(_02030_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07639_ (.I(_02928_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07640_ (.A1(_02930_),
    .A2(_02931_),
    .B(_02923_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07641_ (.A1(_02925_),
    .A2(_02929_),
    .B(_02932_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07642_ (.I(\mem.mem_dff.code_mem[30][1] ),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07643_ (.A1(_02852_),
    .A2(_02931_),
    .B(_02923_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07644_ (.A1(_02933_),
    .A2(_02929_),
    .B(_02934_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07645_ (.I(\mem.mem_dff.code_mem[30][2] ),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07646_ (.I(_02040_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07647_ (.A1(_02936_),
    .A2(_02931_),
    .B(_02923_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07648_ (.A1(_02935_),
    .A2(_02929_),
    .B(_02937_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07649_ (.I(\mem.mem_dff.code_mem[30][3] ),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07650_ (.I(_02897_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07651_ (.A1(_02857_),
    .A2(_02931_),
    .B(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07652_ (.A1(_02938_),
    .A2(_02929_),
    .B(_02940_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07653_ (.I(\mem.mem_dff.code_mem[30][4] ),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07654_ (.I(_02928_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07655_ (.I(_02050_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07656_ (.I(_02928_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07657_ (.A1(_02943_),
    .A2(_02944_),
    .B(_02939_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07658_ (.A1(_02941_),
    .A2(_02942_),
    .B(_02945_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07659_ (.I(\mem.mem_dff.code_mem[30][5] ),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07660_ (.I(_02055_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07661_ (.A1(_02947_),
    .A2(_02944_),
    .B(_02939_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07662_ (.A1(_02946_),
    .A2(_02942_),
    .B(_02948_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07663_ (.I(\mem.mem_dff.code_mem[30][6] ),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07664_ (.A1(_02867_),
    .A2(_02944_),
    .B(_02939_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07665_ (.A1(_02949_),
    .A2(_02942_),
    .B(_02950_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07666_ (.I(\mem.mem_dff.code_mem[30][7] ),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07667_ (.I(_02840_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07668_ (.I(_02952_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07669_ (.A1(_02870_),
    .A2(_02944_),
    .B(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07670_ (.A1(_02951_),
    .A2(_02942_),
    .B(_02954_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07671_ (.I(\mem.mem_dff.code_mem[31][0] ),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07672_ (.A1(_02787_),
    .A2(_02412_),
    .A3(_02255_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07673_ (.I(_02956_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07674_ (.A1(_02874_),
    .A2(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07675_ (.I(_02958_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07676_ (.I(_02958_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07677_ (.A1(_02930_),
    .A2(_02960_),
    .B(_02953_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07678_ (.A1(_02955_),
    .A2(_02959_),
    .B(_02961_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07679_ (.I(\mem.mem_dff.code_mem[31][1] ),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07680_ (.I(_02036_),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07681_ (.A1(_02963_),
    .A2(_02960_),
    .B(_02953_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07682_ (.A1(_02962_),
    .A2(_02959_),
    .B(_02964_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07683_ (.I(\mem.mem_dff.code_mem[31][2] ),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07684_ (.A1(_02936_),
    .A2(_02960_),
    .B(_02953_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07685_ (.A1(_02965_),
    .A2(_02959_),
    .B(_02966_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07686_ (.I(\mem.mem_dff.code_mem[31][3] ),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_02044_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07688_ (.I(_02952_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07689_ (.A1(_02968_),
    .A2(_02960_),
    .B(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07690_ (.A1(_02967_),
    .A2(_02959_),
    .B(_02970_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07691_ (.I(\mem.mem_dff.code_mem[31][4] ),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07692_ (.I(_02958_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07693_ (.I(_02958_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07694_ (.A1(_02943_),
    .A2(_02973_),
    .B(_02969_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07695_ (.A1(_02971_),
    .A2(_02972_),
    .B(_02974_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07696_ (.I(\mem.mem_dff.code_mem[31][5] ),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07697_ (.A1(_02947_),
    .A2(_02973_),
    .B(_02969_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07698_ (.A1(_02975_),
    .A2(_02972_),
    .B(_02976_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07699_ (.I(\mem.mem_dff.code_mem[31][6] ),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07700_ (.I(_02059_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07701_ (.A1(_02978_),
    .A2(_02973_),
    .B(_02969_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07702_ (.A1(_02977_),
    .A2(_02972_),
    .B(_02979_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07703_ (.I(\mem.mem_dff.code_mem[31][7] ),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07704_ (.I(_02063_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07705_ (.I(_02952_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07706_ (.A1(_02981_),
    .A2(_02973_),
    .B(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07707_ (.A1(_02980_),
    .A2(_02972_),
    .B(_02983_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07708_ (.I(_02101_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07709_ (.I(net254),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07710_ (.I(_02021_),
    .Z(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07711_ (.A1(_02345_),
    .A2(net186),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07712_ (.A1(_00764_),
    .A2(_01173_),
    .A3(_01174_),
    .A4(_02987_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07713_ (.A1(_02014_),
    .A2(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07714_ (.A1(_02985_),
    .A2(_02986_),
    .A3(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07715_ (.I(_02990_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07716_ (.I(_02990_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07717_ (.A1(\mem.mem_dff.data_mem[0][0] ),
    .A2(_02992_),
    .B(_02982_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07718_ (.A1(_02984_),
    .A2(_02991_),
    .B(_02993_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07719_ (.I(_02143_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07720_ (.A1(\mem.mem_dff.data_mem[0][1] ),
    .A2(_02992_),
    .B(_02982_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07721_ (.A1(_02994_),
    .A2(_02991_),
    .B(_02995_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07722_ (.I(_02108_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07723_ (.A1(\mem.mem_dff.data_mem[0][2] ),
    .A2(_02992_),
    .B(_02982_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07724_ (.A1(_02996_),
    .A2(_02991_),
    .B(_02997_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07725_ (.I(_02149_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07726_ (.I(_02952_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07727_ (.A1(\mem.mem_dff.data_mem[0][3] ),
    .A2(_02992_),
    .B(_02999_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07728_ (.A1(_02998_),
    .A2(_02991_),
    .B(_03000_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07729_ (.I(_02116_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07730_ (.I(_02990_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07731_ (.I(_02990_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07732_ (.A1(\mem.mem_dff.data_mem[0][4] ),
    .A2(_03003_),
    .B(_02999_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07733_ (.A1(_03001_),
    .A2(_03002_),
    .B(_03004_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07734_ (.I(_02121_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07735_ (.A1(\mem.mem_dff.data_mem[0][5] ),
    .A2(_03003_),
    .B(_02999_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07736_ (.A1(_03005_),
    .A2(_03002_),
    .B(_03006_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07737_ (.I(_02160_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07738_ (.A1(\mem.mem_dff.data_mem[0][6] ),
    .A2(_03003_),
    .B(_02999_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07739_ (.A1(_03007_),
    .A2(_03002_),
    .B(_03008_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07740_ (.I(_02164_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07741_ (.I(_02840_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07742_ (.I(_03010_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07743_ (.A1(\mem.mem_dff.data_mem[0][7] ),
    .A2(_03003_),
    .B(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07744_ (.A1(_03009_),
    .A2(_03002_),
    .B(_03012_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07745_ (.I(\mem.mem_dff.data_mem[1][0] ),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07746_ (.I(_00762_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07747_ (.A1(_02381_),
    .A2(_03014_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07748_ (.I(_03015_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07749_ (.A1(_02014_),
    .A2(_02988_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07750_ (.I(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07751_ (.A1(_03016_),
    .A2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07752_ (.I(_03019_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07753_ (.I(_03019_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07754_ (.A1(_02930_),
    .A2(_03021_),
    .B(_03011_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07755_ (.A1(_03013_),
    .A2(_03020_),
    .B(_03022_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07756_ (.I(\mem.mem_dff.data_mem[1][1] ),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07757_ (.A1(_02963_),
    .A2(_03021_),
    .B(_03011_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07758_ (.A1(_03023_),
    .A2(_03020_),
    .B(_03024_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07759_ (.I(\mem.mem_dff.data_mem[1][2] ),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07760_ (.A1(_02936_),
    .A2(_03021_),
    .B(_03011_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07761_ (.A1(_03025_),
    .A2(_03020_),
    .B(_03026_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07762_ (.I(\mem.mem_dff.data_mem[1][3] ),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07763_ (.I(_03010_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07764_ (.A1(_02968_),
    .A2(_03021_),
    .B(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07765_ (.A1(_03027_),
    .A2(_03020_),
    .B(_03029_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07766_ (.I(\mem.mem_dff.data_mem[1][4] ),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07767_ (.I(_03019_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07768_ (.I(_03019_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07769_ (.A1(_02943_),
    .A2(_03032_),
    .B(_03028_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07770_ (.A1(_03030_),
    .A2(_03031_),
    .B(_03033_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07771_ (.I(\mem.mem_dff.data_mem[1][5] ),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07772_ (.A1(_02947_),
    .A2(_03032_),
    .B(_03028_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07773_ (.A1(_03034_),
    .A2(_03031_),
    .B(_03035_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07774_ (.I(\mem.mem_dff.data_mem[1][6] ),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07775_ (.A1(_02978_),
    .A2(_03032_),
    .B(_03028_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07776_ (.A1(_03036_),
    .A2(_03031_),
    .B(_03037_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07777_ (.I(\mem.mem_dff.data_mem[1][7] ),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07778_ (.I(_03010_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07779_ (.A1(_02981_),
    .A2(_03032_),
    .B(_03039_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07780_ (.A1(_03038_),
    .A2(_03031_),
    .B(_03040_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07781_ (.I(\mem.mem_dff.data_mem[2][0] ),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07782_ (.I(_00761_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07783_ (.A1(_02381_),
    .A2(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07784_ (.I(_03043_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07785_ (.A1(_03044_),
    .A2(_03018_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07786_ (.I(_03045_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07787_ (.I(_03045_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07788_ (.A1(_02930_),
    .A2(_03047_),
    .B(_03039_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07789_ (.A1(_03041_),
    .A2(_03046_),
    .B(_03048_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07790_ (.I(\mem.mem_dff.data_mem[2][1] ),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07791_ (.A1(_02963_),
    .A2(_03047_),
    .B(_03039_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07792_ (.A1(_03049_),
    .A2(_03046_),
    .B(_03050_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07793_ (.I(\mem.mem_dff.data_mem[2][2] ),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07794_ (.A1(_02936_),
    .A2(_03047_),
    .B(_03039_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07795_ (.A1(_03051_),
    .A2(_03046_),
    .B(_03052_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07796_ (.I(\mem.mem_dff.data_mem[2][3] ),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_03010_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07798_ (.A1(_02968_),
    .A2(_03047_),
    .B(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07799_ (.A1(_03053_),
    .A2(_03046_),
    .B(_03055_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07800_ (.I(\mem.mem_dff.data_mem[2][4] ),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07801_ (.I(_03045_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07802_ (.I(_03045_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07803_ (.A1(_02943_),
    .A2(_03058_),
    .B(_03054_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07804_ (.A1(_03056_),
    .A2(_03057_),
    .B(_03059_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07805_ (.I(\mem.mem_dff.data_mem[2][5] ),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07806_ (.A1(_02947_),
    .A2(_03058_),
    .B(_03054_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07807_ (.A1(_03060_),
    .A2(_03057_),
    .B(_03061_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07808_ (.I(\mem.mem_dff.data_mem[2][6] ),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07809_ (.A1(_02978_),
    .A2(_03058_),
    .B(_03054_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07810_ (.A1(_03062_),
    .A2(_03057_),
    .B(_03063_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07811_ (.I(\mem.mem_dff.data_mem[2][7] ),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07812_ (.I(_01998_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07813_ (.I(_03065_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07814_ (.A1(_02981_),
    .A2(_03058_),
    .B(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07815_ (.A1(_03064_),
    .A2(_03057_),
    .B(_03067_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07816_ (.I(\mem.mem_dff.data_mem[3][0] ),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07817_ (.A1(_02381_),
    .A2(_02135_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07818_ (.I(_03069_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(_03070_),
    .A2(_03018_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07820_ (.I(_03071_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07821_ (.I(_02030_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07822_ (.I(_03071_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07823_ (.A1(_03073_),
    .A2(_03074_),
    .B(_03066_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07824_ (.A1(_03068_),
    .A2(_03072_),
    .B(_03075_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07825_ (.I(\mem.mem_dff.data_mem[3][1] ),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07826_ (.A1(_02963_),
    .A2(_03074_),
    .B(_03066_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07827_ (.A1(_03076_),
    .A2(_03072_),
    .B(_03077_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07828_ (.I(\mem.mem_dff.data_mem[3][2] ),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07829_ (.I(_02040_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07830_ (.A1(_03079_),
    .A2(_03074_),
    .B(_03066_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07831_ (.A1(_03078_),
    .A2(_03072_),
    .B(_03080_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07832_ (.I(\mem.mem_dff.data_mem[3][3] ),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07833_ (.I(_03065_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07834_ (.A1(_02968_),
    .A2(_03074_),
    .B(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07835_ (.A1(_03081_),
    .A2(_03072_),
    .B(_03083_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07836_ (.I(\mem.mem_dff.data_mem[3][4] ),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07837_ (.I(_03071_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07838_ (.I(_02050_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07839_ (.I(_03071_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07840_ (.A1(_03086_),
    .A2(_03087_),
    .B(_03082_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07841_ (.A1(_03084_),
    .A2(_03085_),
    .B(_03088_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07842_ (.I(\mem.mem_dff.data_mem[3][5] ),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07843_ (.I(_02055_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07844_ (.A1(_03090_),
    .A2(_03087_),
    .B(_03082_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07845_ (.A1(_03089_),
    .A2(_03085_),
    .B(_03091_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07846_ (.I(\mem.mem_dff.data_mem[3][6] ),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07847_ (.A1(_02978_),
    .A2(_03087_),
    .B(_03082_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07848_ (.A1(_03092_),
    .A2(_03085_),
    .B(_03093_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07849_ (.I(\mem.mem_dff.data_mem[3][7] ),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07850_ (.I(_03065_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07851_ (.A1(_02981_),
    .A2(_03087_),
    .B(_03095_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07852_ (.A1(_03094_),
    .A2(_03085_),
    .B(_03096_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07853_ (.I(\mem.mem_dff.data_mem[4][0] ),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07854_ (.I(_02020_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07855_ (.I(_02289_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07856_ (.A1(_03098_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07857_ (.I(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07858_ (.A1(_03101_),
    .A2(_03018_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07859_ (.I(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07860_ (.I(_03102_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07861_ (.A1(_03073_),
    .A2(_03104_),
    .B(_03095_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07862_ (.A1(_03097_),
    .A2(_03103_),
    .B(_03105_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07863_ (.I(\mem.mem_dff.data_mem[4][1] ),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07864_ (.I(_02036_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07865_ (.A1(_03107_),
    .A2(_03104_),
    .B(_03095_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07866_ (.A1(_03106_),
    .A2(_03103_),
    .B(_03108_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07867_ (.I(\mem.mem_dff.data_mem[4][2] ),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07868_ (.A1(_03079_),
    .A2(_03104_),
    .B(_03095_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07869_ (.A1(_03109_),
    .A2(_03103_),
    .B(_03110_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07870_ (.I(\mem.mem_dff.data_mem[4][3] ),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07871_ (.I(_02044_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07872_ (.I(_03065_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07873_ (.A1(_03112_),
    .A2(_03104_),
    .B(_03113_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07874_ (.A1(_03111_),
    .A2(_03103_),
    .B(_03114_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07875_ (.I(\mem.mem_dff.data_mem[4][4] ),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07876_ (.I(_03102_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07877_ (.I(_03102_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07878_ (.A1(_03086_),
    .A2(_03117_),
    .B(_03113_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07879_ (.A1(_03115_),
    .A2(_03116_),
    .B(_03118_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07880_ (.I(\mem.mem_dff.data_mem[4][5] ),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07881_ (.A1(_03090_),
    .A2(_03117_),
    .B(_03113_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07882_ (.A1(_03119_),
    .A2(_03116_),
    .B(_03120_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07883_ (.I(\mem.mem_dff.data_mem[4][6] ),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07884_ (.I(_02059_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07885_ (.A1(_03122_),
    .A2(_03117_),
    .B(_03113_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07886_ (.A1(_03121_),
    .A2(_03116_),
    .B(_03123_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07887_ (.I(\mem.mem_dff.data_mem[4][7] ),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07888_ (.I(_02063_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07889_ (.I(_01998_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07890_ (.I(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07891_ (.A1(_03125_),
    .A2(_03117_),
    .B(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07892_ (.A1(_03124_),
    .A2(_03116_),
    .B(_03128_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07893_ (.I(\mem.mem_dff.data_mem[5][0] ),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07894_ (.A1(_02020_),
    .A2(_03014_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07895_ (.I(_03130_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07896_ (.A1(_03131_),
    .A2(_03017_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07897_ (.I(_03132_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07898_ (.I(_03132_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07899_ (.A1(_03073_),
    .A2(_03134_),
    .B(_03127_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07900_ (.A1(_03129_),
    .A2(_03133_),
    .B(_03135_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07901_ (.I(\mem.mem_dff.data_mem[5][1] ),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07902_ (.A1(_03107_),
    .A2(_03134_),
    .B(_03127_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07903_ (.A1(_03136_),
    .A2(_03133_),
    .B(_03137_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07904_ (.I(\mem.mem_dff.data_mem[5][2] ),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07905_ (.A1(_03079_),
    .A2(_03134_),
    .B(_03127_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07906_ (.A1(_03138_),
    .A2(_03133_),
    .B(_03139_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07907_ (.I(\mem.mem_dff.data_mem[5][3] ),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07908_ (.I(_03126_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07909_ (.A1(_03112_),
    .A2(_03134_),
    .B(_03141_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07910_ (.A1(_03140_),
    .A2(_03133_),
    .B(_03142_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07911_ (.I(\mem.mem_dff.data_mem[5][4] ),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07912_ (.I(_03132_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07913_ (.I(_03132_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07914_ (.A1(_03086_),
    .A2(_03145_),
    .B(_03141_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07915_ (.A1(_03143_),
    .A2(_03144_),
    .B(_03146_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07916_ (.I(\mem.mem_dff.data_mem[5][5] ),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07917_ (.A1(_03090_),
    .A2(_03145_),
    .B(_03141_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07918_ (.A1(_03147_),
    .A2(_03144_),
    .B(_03148_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07919_ (.I(\mem.mem_dff.data_mem[5][6] ),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07920_ (.A1(_03122_),
    .A2(_03145_),
    .B(_03141_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07921_ (.A1(_03149_),
    .A2(_03144_),
    .B(_03150_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07922_ (.I(\mem.mem_dff.data_mem[5][7] ),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07923_ (.I(_03126_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07924_ (.A1(_03125_),
    .A2(_03145_),
    .B(_03152_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07925_ (.A1(_03151_),
    .A2(_03144_),
    .B(_03153_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07926_ (.A1(_02467_),
    .A2(_02989_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07927_ (.I(_03154_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07928_ (.I(_03154_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07929_ (.A1(\mem.mem_dff.data_mem[6][0] ),
    .A2(_03156_),
    .B(_03152_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07930_ (.A1(_02984_),
    .A2(_03155_),
    .B(_03157_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07931_ (.A1(\mem.mem_dff.data_mem[6][1] ),
    .A2(_03156_),
    .B(_03152_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07932_ (.A1(_02994_),
    .A2(_03155_),
    .B(_03158_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07933_ (.A1(\mem.mem_dff.data_mem[6][2] ),
    .A2(_03156_),
    .B(_03152_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07934_ (.A1(_02996_),
    .A2(_03155_),
    .B(_03159_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07935_ (.I(_03126_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07936_ (.A1(\mem.mem_dff.data_mem[6][3] ),
    .A2(_03156_),
    .B(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07937_ (.A1(_02998_),
    .A2(_03155_),
    .B(_03161_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07938_ (.I(_03154_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07939_ (.I(_03154_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07940_ (.A1(\mem.mem_dff.data_mem[6][4] ),
    .A2(_03163_),
    .B(_03160_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07941_ (.A1(_03001_),
    .A2(_03162_),
    .B(_03164_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07942_ (.A1(\mem.mem_dff.data_mem[6][5] ),
    .A2(_03163_),
    .B(_03160_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07943_ (.A1(_03005_),
    .A2(_03162_),
    .B(_03165_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07944_ (.A1(\mem.mem_dff.data_mem[6][6] ),
    .A2(_03163_),
    .B(_03160_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07945_ (.A1(_03007_),
    .A2(_03162_),
    .B(_03166_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07946_ (.I(_01998_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07947_ (.I(_03167_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07948_ (.A1(\mem.mem_dff.data_mem[6][7] ),
    .A2(_03163_),
    .B(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07949_ (.A1(_03009_),
    .A2(_03162_),
    .B(_03169_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07950_ (.A1(_02256_),
    .A2(_02989_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07951_ (.I(_03170_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07952_ (.I(_03170_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07953_ (.A1(\mem.mem_dff.data_mem[7][0] ),
    .A2(_03172_),
    .B(_03168_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07954_ (.A1(_02984_),
    .A2(_03171_),
    .B(_03173_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07955_ (.A1(\mem.mem_dff.data_mem[7][1] ),
    .A2(_03172_),
    .B(_03168_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07956_ (.A1(_02994_),
    .A2(_03171_),
    .B(_03174_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07957_ (.A1(\mem.mem_dff.data_mem[7][2] ),
    .A2(_03172_),
    .B(_03168_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07958_ (.A1(_02996_),
    .A2(_03171_),
    .B(_03175_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07959_ (.I(_03167_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07960_ (.A1(\mem.mem_dff.data_mem[7][3] ),
    .A2(_03172_),
    .B(_03176_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07961_ (.A1(_02998_),
    .A2(_03171_),
    .B(_03177_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07962_ (.I(_03170_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07963_ (.I(_03170_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07964_ (.A1(\mem.mem_dff.data_mem[7][4] ),
    .A2(_03179_),
    .B(_03176_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07965_ (.A1(_03001_),
    .A2(_03178_),
    .B(_03180_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07966_ (.A1(\mem.mem_dff.data_mem[7][5] ),
    .A2(_03179_),
    .B(_03176_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07967_ (.A1(_03005_),
    .A2(_03178_),
    .B(_03181_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07968_ (.A1(\mem.mem_dff.data_mem[7][6] ),
    .A2(_03179_),
    .B(_03176_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07969_ (.A1(_03007_),
    .A2(_03178_),
    .B(_03182_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07970_ (.I(_03167_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07971_ (.A1(\mem.mem_dff.data_mem[7][7] ),
    .A2(_03179_),
    .B(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07972_ (.A1(_03009_),
    .A2(_03178_),
    .B(_03184_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07973_ (.I(_02002_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07974_ (.I(_01675_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07975_ (.I(_01683_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07976_ (.I(_03187_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07977_ (.I(_01691_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07978_ (.A1(_01699_),
    .A2(_01703_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07979_ (.I(_01710_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07980_ (.A1(_03190_),
    .A2(_03191_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07981_ (.A1(_03186_),
    .A2(_03188_),
    .A3(_03189_),
    .A4(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07982_ (.I(_01605_),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07983_ (.I(_01616_),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07984_ (.A1(_01597_),
    .A2(_01606_),
    .A3(_01615_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07985_ (.A1(_01587_),
    .A2(_03196_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07986_ (.A1(_03194_),
    .A2(_03195_),
    .A3(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07987_ (.I(_01701_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07988_ (.A1(_01633_),
    .A2(_01635_),
    .A3(_01604_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07989_ (.A1(_03199_),
    .A2(_03200_),
    .Z(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07990_ (.I(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07991_ (.A1(_03198_),
    .A2(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07992_ (.A1(_03185_),
    .A2(_03193_),
    .A3(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07993_ (.I(_03204_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07994_ (.A1(\stack[28][0] ),
    .A2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07995_ (.I(_01756_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07996_ (.I(_03207_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07997_ (.I(_03193_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07998_ (.I(_03203_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07999_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03210_),
    .B2(net144),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08000_ (.A1(_03206_),
    .A2(_03211_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08001_ (.I(_03210_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08002_ (.I(_03212_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08003_ (.I(_01791_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08004_ (.I(_03214_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08005_ (.A1(_03215_),
    .A2(_03209_),
    .B1(_03205_),
    .B2(\stack[28][1] ),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08006_ (.A1(_01764_),
    .A2(_03213_),
    .B(_03216_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08007_ (.I(_01823_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08008_ (.I(_03217_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08009_ (.A1(_03218_),
    .A2(_03209_),
    .B1(_03205_),
    .B2(\stack[28][2] ),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08010_ (.A1(_01797_),
    .A2(_03213_),
    .B(_03219_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08011_ (.I(_01855_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08012_ (.I(_03220_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08013_ (.A1(_03221_),
    .A2(_03209_),
    .B1(_03205_),
    .B2(\stack[28][3] ),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08014_ (.A1(_01829_),
    .A2(_03213_),
    .B(_03222_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08015_ (.I(_01886_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08016_ (.I(_03223_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08017_ (.I(_03204_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08018_ (.A1(_03224_),
    .A2(_03193_),
    .B1(_03225_),
    .B2(\stack[28][4] ),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08019_ (.A1(_01861_),
    .A2(_03213_),
    .B(_03226_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08020_ (.I(_01921_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08021_ (.I(_03227_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08022_ (.A1(_03228_),
    .A2(_03193_),
    .B1(_03225_),
    .B2(\stack[28][5] ),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08023_ (.A1(_01893_),
    .A2(_03212_),
    .B(_03229_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08024_ (.I(_01692_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08025_ (.A1(_01677_),
    .A2(_01925_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08026_ (.A1(_03230_),
    .A2(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08027_ (.A1(_03190_),
    .A2(_01711_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08028_ (.I(_03233_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08029_ (.I(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08030_ (.A1(_03232_),
    .A2(_03235_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08031_ (.I(_01123_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08032_ (.I(_03237_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08033_ (.A1(_03238_),
    .A2(_03210_),
    .B1(_03225_),
    .B2(\stack[28][6] ),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08034_ (.A1(_01964_),
    .A2(_03236_),
    .B(_03239_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08035_ (.A1(net152),
    .A2(_03210_),
    .B1(_03225_),
    .B2(\stack[28][7] ),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08036_ (.A1(_01991_),
    .A2(_03236_),
    .B(_03240_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(_00763_),
    .A2(_01177_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08038_ (.I(_03241_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08039_ (.I(_03242_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08040_ (.I(_03243_),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08041_ (.A1(net253),
    .A2(_03243_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08042_ (.I(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08043_ (.A1(_02345_),
    .A2(net188),
    .A3(_01174_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08044_ (.I(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08045_ (.A1(_02985_),
    .A2(_02256_),
    .A3(_03248_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08046_ (.I(_03249_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08047_ (.A1(_02985_),
    .A2(_02467_),
    .A3(_03248_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08048_ (.I(_03251_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08049_ (.A1(_02291_),
    .A2(_03248_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08050_ (.I(_03253_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08051_ (.A1(net69),
    .A2(_03252_),
    .B1(_03254_),
    .B2(net120),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08052_ (.A1(net112),
    .A2(_03250_),
    .B(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08053_ (.A1(\mem.io_data_out[0] ),
    .A2(_03244_),
    .B1(_03246_),
    .B2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08054_ (.A1(_02005_),
    .A2(_03257_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08055_ (.A1(net70),
    .A2(_03252_),
    .B1(_03254_),
    .B2(net121),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08056_ (.A1(net113),
    .A2(_03250_),
    .B(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08057_ (.A1(\mem.io_data_out[1] ),
    .A2(_03244_),
    .B1(_03246_),
    .B2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08058_ (.A1(_02005_),
    .A2(_03260_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08059_ (.I(_02002_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08060_ (.I(_03261_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08061_ (.I(_03262_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08062_ (.A1(net71),
    .A2(_03252_),
    .B1(_03254_),
    .B2(net122),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08063_ (.A1(net114),
    .A2(_03250_),
    .B(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08064_ (.A1(\mem.io_data_out[2] ),
    .A2(_03244_),
    .B1(_03246_),
    .B2(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08065_ (.A1(_03263_),
    .A2(_03266_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08066_ (.I(_03243_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08067_ (.A1(net72),
    .A2(_03252_),
    .B1(_03254_),
    .B2(net123),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08068_ (.A1(net115),
    .A2(_03250_),
    .B(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08069_ (.A1(\mem.io_data_out[3] ),
    .A2(_03267_),
    .B1(_03246_),
    .B2(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08070_ (.A1(_03263_),
    .A2(_03270_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08071_ (.I(_03245_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(_03249_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08073_ (.I(_03251_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08074_ (.I(_03253_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08075_ (.A1(net73),
    .A2(_03273_),
    .B1(_03274_),
    .B2(net124),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08076_ (.A1(net116),
    .A2(_03272_),
    .B(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08077_ (.A1(\mem.io_data_out[4] ),
    .A2(_03267_),
    .B1(_03271_),
    .B2(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08078_ (.A1(_03263_),
    .A2(_03277_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08079_ (.A1(net74),
    .A2(_03273_),
    .B1(_03274_),
    .B2(net125),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08080_ (.A1(net117),
    .A2(_03272_),
    .B(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08081_ (.A1(\mem.io_data_out[5] ),
    .A2(_03267_),
    .B1(_03271_),
    .B2(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08082_ (.A1(_03263_),
    .A2(_03280_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08083_ (.I(_03261_),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08084_ (.I(_03281_),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08085_ (.A1(net75),
    .A2(_03273_),
    .B1(_03274_),
    .B2(net126),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08086_ (.A1(net118),
    .A2(_03272_),
    .B(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08087_ (.A1(\mem.io_data_out[6] ),
    .A2(_03267_),
    .B1(_03271_),
    .B2(_03284_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08088_ (.A1(_03282_),
    .A2(_03285_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08089_ (.A1(net76),
    .A2(_03273_),
    .B1(_03274_),
    .B2(net127),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08090_ (.A1(net119),
    .A2(_03272_),
    .B(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08091_ (.A1(\mem.io_data_out[7] ),
    .A2(_03243_),
    .B1(_03271_),
    .B2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08092_ (.A1(_03282_),
    .A2(_03288_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08093_ (.A1(_02290_),
    .A2(_02987_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08094_ (.I(_03289_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(\mem.mem_dff.code_mem[23][0] ),
    .A2(_02731_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08096_ (.I(_02292_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08097_ (.I(_02700_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08098_ (.A1(\mem.mem_dff.code_mem[8][0] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\mem.mem_dff.code_mem[22][0] ),
    .C1(\mem.mem_dff.code_mem[31][0] ),
    .C2(_02957_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08099_ (.A1(\mem.mem_dff.code_mem[15][0] ),
    .A2(_02499_),
    .B1(_02902_),
    .B2(\mem.mem_dff.code_mem[29][0] ),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08100_ (.A1(\mem.mem_dff.code_mem[6][0] ),
    .A2(_02226_),
    .B1(_02927_),
    .B2(\mem.mem_dff.code_mem[30][0] ),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08101_ (.A1(_03291_),
    .A2(_03294_),
    .A3(_03295_),
    .A4(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08102_ (.A1(\mem.mem_dff.code_mem[9][0] ),
    .A2(_02321_),
    .B1(_02876_),
    .B2(\mem.mem_dff.code_mem[28][0] ),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08103_ (.I(_02382_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08104_ (.I(_02814_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08105_ (.A1(\mem.mem_dff.code_mem[12][0] ),
    .A2(_02413_),
    .B1(_02441_),
    .B2(\mem.mem_dff.code_mem[13][0] ),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08106_ (.A1(\mem.mem_dff.code_mem[10][0] ),
    .A2(_02346_),
    .B1(_02761_),
    .B2(\mem.mem_dff.code_mem[24][0] ),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08107_ (.A1(\mem.mem_dff.code_mem[25][0] ),
    .A2(_02788_),
    .B1(_02845_),
    .B2(\mem.mem_dff.code_mem[27][0] ),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08108_ (.A1(_03301_),
    .A2(_03302_),
    .A3(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08109_ (.A1(\mem.mem_dff.code_mem[11][0] ),
    .A2(_03299_),
    .B1(_03300_),
    .B2(\mem.mem_dff.code_mem[26][0] ),
    .C(_03304_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08110_ (.A1(\mem.mem_dff.code_mem[1][0] ),
    .A2(_02070_),
    .B1(_02561_),
    .B2(\mem.mem_dff.code_mem[17][0] ),
    .C(_02026_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08111_ (.I(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08112_ (.A1(\mem.mem_dff.code_mem[5][0] ),
    .A2(_02199_),
    .B1(_02649_),
    .B2(\mem.mem_dff.code_mem[20][0] ),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08113_ (.A1(\mem.mem_dff.code_mem[2][0] ),
    .A2(_02097_),
    .B1(_02587_),
    .B2(\mem.mem_dff.code_mem[18][0] ),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08114_ (.A1(\mem.mem_dff.code_mem[19][0] ),
    .A2(_02619_),
    .B1(_02675_),
    .B2(\mem.mem_dff.code_mem[21][0] ),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08115_ (.A1(\mem.mem_dff.code_mem[3][0] ),
    .A2(_02136_),
    .B1(_02172_),
    .B2(\mem.mem_dff.code_mem[4][0] ),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08116_ (.A1(_03308_),
    .A2(_03309_),
    .A3(_03310_),
    .A4(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08117_ (.A1(\mem.mem_dff.code_mem[16][0] ),
    .A2(_02536_),
    .B(_03307_),
    .C(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08118_ (.A1(\mem.mem_dff.code_mem[7][0] ),
    .A2(_02258_),
    .B1(_02469_),
    .B2(\mem.mem_dff.code_mem[14][0] ),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08119_ (.A1(_03298_),
    .A2(_03305_),
    .A3(_03313_),
    .A4(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08120_ (.I(_02015_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08121_ (.A1(\mem.mem_dff.code_mem[0][0] ),
    .A2(_03290_),
    .B1(_03297_),
    .B2(_03315_),
    .C(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08122_ (.I(_02986_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08123_ (.I(_02988_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08124_ (.A1(_03098_),
    .A2(_02135_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08125_ (.I(_03320_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08126_ (.A1(\mem.mem_dff.data_mem[1][0] ),
    .A2(_03016_),
    .B1(_03070_),
    .B2(\mem.mem_dff.data_mem[3][0] ),
    .C1(\mem.mem_dff.data_mem[7][0] ),
    .C2(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08127_ (.I(_03100_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08128_ (.I(_03130_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08129_ (.I(_02290_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08130_ (.A1(\mem.mem_dff.data_mem[4][0] ),
    .A2(_03323_),
    .B1(_03324_),
    .B2(\mem.mem_dff.data_mem[5][0] ),
    .C(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08131_ (.I(_03043_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08132_ (.A1(_03098_),
    .A2(_03042_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08133_ (.I(_03328_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08134_ (.A1(\mem.mem_dff.data_mem[2][0] ),
    .A2(_03327_),
    .B1(_03329_),
    .B2(\mem.mem_dff.data_mem[6][0] ),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08135_ (.A1(_03322_),
    .A2(_03326_),
    .A3(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08136_ (.A1(\mem.mem_dff.data_mem[0][0] ),
    .A2(_03318_),
    .B(_03319_),
    .C(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(_03317_),
    .A2(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08138_ (.A1(_01995_),
    .A2(_01996_),
    .B(_02008_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08139_ (.A1(_02014_),
    .A2(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08140_ (.I(_03335_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08141_ (.I0(\mem.dff_data_out[0] ),
    .I1(_03333_),
    .S(_03336_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08142_ (.I(_03337_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08143_ (.A1(\mem.mem_dff.code_mem[9][1] ),
    .A2(_02321_),
    .B1(_02876_),
    .B2(\mem.mem_dff.code_mem[28][1] ),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08144_ (.A1(\mem.mem_dff.code_mem[7][1] ),
    .A2(_02258_),
    .B1(_02469_),
    .B2(\mem.mem_dff.code_mem[14][1] ),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08145_ (.I(_02788_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08146_ (.I(_02845_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08147_ (.A1(\mem.mem_dff.code_mem[25][1] ),
    .A2(_03340_),
    .B1(_03341_),
    .B2(\mem.mem_dff.code_mem[27][1] ),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08148_ (.I(_02346_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08149_ (.I(_02761_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08150_ (.A1(\mem.mem_dff.code_mem[10][1] ),
    .A2(_03343_),
    .B1(_03344_),
    .B2(\mem.mem_dff.code_mem[24][1] ),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08151_ (.A1(\mem.mem_dff.code_mem[12][1] ),
    .A2(_02414_),
    .B1(_02442_),
    .B2(\mem.mem_dff.code_mem[13][1] ),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08152_ (.A1(_03342_),
    .A2(_03345_),
    .A3(_03346_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08153_ (.A1(\mem.mem_dff.code_mem[11][1] ),
    .A2(_02383_),
    .B1(_02815_),
    .B2(\mem.mem_dff.code_mem[26][1] ),
    .C(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08154_ (.I(_02097_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08155_ (.I(_02587_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08156_ (.A1(\mem.mem_dff.code_mem[2][1] ),
    .A2(_03349_),
    .B1(_03350_),
    .B2(\mem.mem_dff.code_mem[18][1] ),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08157_ (.I(_02199_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08158_ (.I(_02649_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08159_ (.A1(\mem.mem_dff.code_mem[5][1] ),
    .A2(_03352_),
    .B1(_03353_),
    .B2(\mem.mem_dff.code_mem[20][1] ),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08160_ (.I(_02070_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08161_ (.I(_02026_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08162_ (.A1(\mem.mem_dff.code_mem[1][1] ),
    .A2(_03355_),
    .B1(_02535_),
    .B2(\mem.mem_dff.code_mem[16][1] ),
    .C(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08163_ (.I(_02561_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08164_ (.I(_02675_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08165_ (.A1(\mem.mem_dff.code_mem[17][1] ),
    .A2(_03358_),
    .B1(_03359_),
    .B2(\mem.mem_dff.code_mem[21][1] ),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08166_ (.A1(_03351_),
    .A2(_03354_),
    .A3(_03357_),
    .A4(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08167_ (.A1(\mem.mem_dff.code_mem[8][1] ),
    .A2(_02292_),
    .B1(_02700_),
    .B2(\mem.mem_dff.code_mem[22][1] ),
    .C1(\mem.mem_dff.code_mem[31][1] ),
    .C2(_02957_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08168_ (.A1(\mem.mem_dff.code_mem[6][1] ),
    .A2(_02226_),
    .B1(_02731_),
    .B2(\mem.mem_dff.code_mem[23][1] ),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02136_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08170_ (.I(_02172_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08171_ (.I(_02619_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08172_ (.A1(\mem.mem_dff.code_mem[3][1] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\mem.mem_dff.code_mem[4][1] ),
    .C1(\mem.mem_dff.code_mem[19][1] ),
    .C2(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08173_ (.I(_02498_),
    .Z(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08174_ (.I(_02901_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08175_ (.A1(\mem.mem_dff.code_mem[15][1] ),
    .A2(_03368_),
    .B1(_03369_),
    .B2(\mem.mem_dff.code_mem[29][1] ),
    .C1(\mem.mem_dff.code_mem[30][1] ),
    .C2(_02927_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08176_ (.A1(_03362_),
    .A2(_03363_),
    .A3(_03367_),
    .A4(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08177_ (.A1(_03361_),
    .A2(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08178_ (.A1(_03338_),
    .A2(_03339_),
    .A3(_03348_),
    .A4(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08179_ (.A1(\mem.mem_dff.code_mem[0][1] ),
    .A2(_03290_),
    .B(_03373_),
    .C(_03316_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08180_ (.I(_03328_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08181_ (.A1(\mem.mem_dff.data_mem[2][1] ),
    .A2(_03044_),
    .B1(_03375_),
    .B2(\mem.mem_dff.data_mem[6][1] ),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08182_ (.I(_03015_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08183_ (.I(_03069_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08184_ (.I(_03320_),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08185_ (.A1(\mem.mem_dff.data_mem[1][1] ),
    .A2(_03377_),
    .B1(_03378_),
    .B2(\mem.mem_dff.data_mem[3][1] ),
    .C1(\mem.mem_dff.data_mem[7][1] ),
    .C2(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08186_ (.I(_02290_),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08187_ (.A1(\mem.mem_dff.data_mem[4][1] ),
    .A2(_03101_),
    .B1(_03131_),
    .B2(\mem.mem_dff.data_mem[5][1] ),
    .C(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08188_ (.A1(_03376_),
    .A2(_03380_),
    .A3(_03382_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08189_ (.A1(\mem.mem_dff.data_mem[0][1] ),
    .A2(_03318_),
    .B(_03319_),
    .C(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08190_ (.A1(_03374_),
    .A2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08191_ (.I0(\mem.dff_data_out[1] ),
    .I1(_03385_),
    .S(_03336_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08192_ (.I(_03386_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08193_ (.A1(\mem.mem_dff.code_mem[15][2] ),
    .A2(_02499_),
    .B1(_02902_),
    .B2(\mem.mem_dff.code_mem[29][2] ),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08194_ (.I(_02225_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08195_ (.I(_02926_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08196_ (.A1(\mem.mem_dff.code_mem[6][2] ),
    .A2(_03388_),
    .B1(_03389_),
    .B2(\mem.mem_dff.code_mem[30][2] ),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08197_ (.I(_02730_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08198_ (.I(_02956_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08199_ (.A1(\mem.mem_dff.code_mem[23][2] ),
    .A2(_03391_),
    .B1(_03392_),
    .B2(\mem.mem_dff.code_mem[31][2] ),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08200_ (.A1(_03387_),
    .A2(_03390_),
    .A3(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08201_ (.A1(\mem.mem_dff.code_mem[8][2] ),
    .A2(_02293_),
    .B1(_02701_),
    .B2(\mem.mem_dff.code_mem[22][2] ),
    .C(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08202_ (.A1(\mem.mem_dff.code_mem[10][2] ),
    .A2(_02347_),
    .B1(_02762_),
    .B2(\mem.mem_dff.code_mem[24][2] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08203_ (.A1(\mem.mem_dff.code_mem[25][2] ),
    .A2(_03340_),
    .B1(_03341_),
    .B2(\mem.mem_dff.code_mem[27][2] ),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08204_ (.A1(\mem.mem_dff.code_mem[12][2] ),
    .A2(_02414_),
    .B1(_02442_),
    .B2(\mem.mem_dff.code_mem[13][2] ),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08205_ (.A1(_03396_),
    .A2(_03397_),
    .A3(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08206_ (.A1(\mem.mem_dff.code_mem[11][2] ),
    .A2(_02383_),
    .B1(_02815_),
    .B2(\mem.mem_dff.code_mem[26][2] ),
    .C(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(_03395_),
    .A2(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08208_ (.A1(\mem.mem_dff.code_mem[3][2] ),
    .A2(_02137_),
    .B1(_02173_),
    .B2(\mem.mem_dff.code_mem[4][2] ),
    .C1(\mem.mem_dff.code_mem[21][2] ),
    .C2(_02676_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08209_ (.A1(\mem.mem_dff.code_mem[5][2] ),
    .A2(_02200_),
    .B1(_02650_),
    .B2(\mem.mem_dff.code_mem[20][2] ),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08210_ (.A1(\mem.mem_dff.code_mem[2][2] ),
    .A2(_02098_),
    .B1(_02588_),
    .B2(\mem.mem_dff.code_mem[18][2] ),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08211_ (.I(_02535_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08212_ (.A1(\mem.mem_dff.code_mem[1][2] ),
    .A2(_03355_),
    .B1(_03405_),
    .B2(\mem.mem_dff.code_mem[16][2] ),
    .C(_03356_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08213_ (.A1(\mem.mem_dff.code_mem[17][2] ),
    .A2(_03358_),
    .B1(_02620_),
    .B2(\mem.mem_dff.code_mem[19][2] ),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08214_ (.A1(_03403_),
    .A2(_03404_),
    .A3(_03406_),
    .A4(_03407_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08215_ (.A1(\mem.mem_dff.code_mem[9][2] ),
    .A2(_02321_),
    .B1(_02876_),
    .B2(\mem.mem_dff.code_mem[28][2] ),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08216_ (.A1(\mem.mem_dff.code_mem[7][2] ),
    .A2(_02258_),
    .B1(_02469_),
    .B2(\mem.mem_dff.code_mem[14][2] ),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08217_ (.A1(_03402_),
    .A2(_03408_),
    .A3(_03409_),
    .A4(_03410_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08218_ (.A1(\mem.mem_dff.code_mem[0][2] ),
    .A2(_03290_),
    .B1(_03401_),
    .B2(_03411_),
    .C(_03316_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08219_ (.A1(\mem.mem_dff.data_mem[2][2] ),
    .A2(_03044_),
    .B1(_03375_),
    .B2(\mem.mem_dff.data_mem[6][2] ),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08220_ (.A1(\mem.mem_dff.data_mem[1][2] ),
    .A2(_03377_),
    .B1(_03378_),
    .B2(\mem.mem_dff.data_mem[3][2] ),
    .C1(\mem.mem_dff.data_mem[7][2] ),
    .C2(_03379_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08221_ (.A1(\mem.mem_dff.data_mem[4][2] ),
    .A2(_03101_),
    .B1(_03131_),
    .B2(\mem.mem_dff.data_mem[5][2] ),
    .C(_03381_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08222_ (.A1(_03413_),
    .A2(_03414_),
    .A3(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08223_ (.A1(\mem.mem_dff.data_mem[0][2] ),
    .A2(_03318_),
    .B(_03319_),
    .C(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(_03412_),
    .A2(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08225_ (.I0(\mem.dff_data_out[2] ),
    .I1(_03418_),
    .S(_03336_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08226_ (.I(_03419_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08227_ (.A1(\mem.mem_dff.code_mem[15][3] ),
    .A2(_03368_),
    .B1(_03369_),
    .B2(\mem.mem_dff.code_mem[29][3] ),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08228_ (.A1(\mem.mem_dff.code_mem[6][3] ),
    .A2(_03388_),
    .B1(_03389_),
    .B2(\mem.mem_dff.code_mem[30][3] ),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08229_ (.A1(\mem.mem_dff.code_mem[23][3] ),
    .A2(_03391_),
    .B1(_03392_),
    .B2(\mem.mem_dff.code_mem[31][3] ),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08230_ (.A1(_03420_),
    .A2(_03421_),
    .A3(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08231_ (.A1(\mem.mem_dff.code_mem[8][3] ),
    .A2(_02293_),
    .B1(_02701_),
    .B2(\mem.mem_dff.code_mem[22][3] ),
    .C(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08232_ (.A1(\mem.mem_dff.code_mem[10][3] ),
    .A2(_02347_),
    .B1(_02762_),
    .B2(\mem.mem_dff.code_mem[24][3] ),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08233_ (.I(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08234_ (.A1(\mem.mem_dff.code_mem[25][3] ),
    .A2(_02789_),
    .B1(_02846_),
    .B2(\mem.mem_dff.code_mem[27][3] ),
    .C(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08235_ (.I(_02257_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08236_ (.I(_02320_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08237_ (.I(_02875_),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08238_ (.A1(\mem.mem_dff.code_mem[7][3] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\mem.mem_dff.code_mem[9][3] ),
    .C1(\mem.mem_dff.code_mem[28][3] ),
    .C2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08239_ (.I(_02468_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08240_ (.A1(\mem.mem_dff.code_mem[12][3] ),
    .A2(_02415_),
    .B1(_03432_),
    .B2(\mem.mem_dff.code_mem[14][3] ),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08241_ (.A1(_03424_),
    .A2(_03427_),
    .A3(_03431_),
    .A4(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08242_ (.A1(\mem.mem_dff.code_mem[3][3] ),
    .A2(_02137_),
    .B1(_02173_),
    .B2(\mem.mem_dff.code_mem[4][3] ),
    .C1(\mem.mem_dff.code_mem[21][3] ),
    .C2(_02676_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08243_ (.A1(\mem.mem_dff.code_mem[5][3] ),
    .A2(_02200_),
    .B1(_02650_),
    .B2(\mem.mem_dff.code_mem[20][3] ),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08244_ (.A1(\mem.mem_dff.code_mem[2][3] ),
    .A2(_02098_),
    .B1(_02588_),
    .B2(\mem.mem_dff.code_mem[18][3] ),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08245_ (.A1(\mem.mem_dff.code_mem[1][3] ),
    .A2(_02071_),
    .B1(_03405_),
    .B2(\mem.mem_dff.code_mem[16][3] ),
    .C(_02027_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08246_ (.A1(\mem.mem_dff.code_mem[17][3] ),
    .A2(_02562_),
    .B1(_02620_),
    .B2(\mem.mem_dff.code_mem[19][3] ),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08247_ (.A1(_03436_),
    .A2(_03437_),
    .A3(_03438_),
    .A4(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _08248_ (.A1(\mem.mem_dff.code_mem[11][3] ),
    .A2(_03299_),
    .B1(_02443_),
    .B2(\mem.mem_dff.code_mem[13][3] ),
    .C1(\mem.mem_dff.code_mem[26][3] ),
    .C2(_03300_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08249_ (.A1(_03435_),
    .A2(_03440_),
    .A3(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08250_ (.A1(\mem.mem_dff.code_mem[0][3] ),
    .A2(_03290_),
    .B1(_03434_),
    .B2(_03442_),
    .C(_03316_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08251_ (.A1(\mem.mem_dff.data_mem[2][3] ),
    .A2(_03044_),
    .B1(_03375_),
    .B2(\mem.mem_dff.data_mem[6][3] ),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08252_ (.A1(\mem.mem_dff.data_mem[1][3] ),
    .A2(_03377_),
    .B1(_03378_),
    .B2(\mem.mem_dff.data_mem[3][3] ),
    .C1(\mem.mem_dff.data_mem[7][3] ),
    .C2(_03379_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08253_ (.A1(\mem.mem_dff.data_mem[4][3] ),
    .A2(_03101_),
    .B1(_03131_),
    .B2(\mem.mem_dff.data_mem[5][3] ),
    .C(_03381_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08254_ (.A1(_03444_),
    .A2(_03445_),
    .A3(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08255_ (.A1(\mem.mem_dff.data_mem[0][3] ),
    .A2(_03318_),
    .B(_03319_),
    .C(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(_03443_),
    .A2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08257_ (.I0(\mem.dff_data_out[3] ),
    .I1(_03449_),
    .S(_03336_),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08258_ (.I(_03450_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08259_ (.I(_03289_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08260_ (.A1(\mem.mem_dff.code_mem[23][4] ),
    .A2(_02731_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08261_ (.A1(\mem.mem_dff.code_mem[8][4] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\mem.mem_dff.code_mem[22][4] ),
    .C1(\mem.mem_dff.code_mem[31][4] ),
    .C2(_02957_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08262_ (.A1(\mem.mem_dff.code_mem[15][4] ),
    .A2(_02499_),
    .B1(_02902_),
    .B2(\mem.mem_dff.code_mem[29][4] ),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08263_ (.A1(\mem.mem_dff.code_mem[6][4] ),
    .A2(_02226_),
    .B1(_02927_),
    .B2(\mem.mem_dff.code_mem[30][4] ),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08264_ (.A1(_03452_),
    .A2(_03453_),
    .A3(_03454_),
    .A4(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08265_ (.A1(\mem.mem_dff.code_mem[10][4] ),
    .A2(_02347_),
    .B1(_02762_),
    .B2(\mem.mem_dff.code_mem[24][4] ),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08266_ (.A1(\mem.mem_dff.code_mem[25][4] ),
    .A2(_03340_),
    .B1(_03341_),
    .B2(\mem.mem_dff.code_mem[27][4] ),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08267_ (.A1(\mem.mem_dff.code_mem[12][4] ),
    .A2(_02413_),
    .B1(_02441_),
    .B2(\mem.mem_dff.code_mem[13][4] ),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08268_ (.A1(_03457_),
    .A2(_03458_),
    .A3(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08269_ (.A1(\mem.mem_dff.code_mem[11][4] ),
    .A2(_02383_),
    .B1(_02815_),
    .B2(\mem.mem_dff.code_mem[26][4] ),
    .C(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08270_ (.A1(\mem.mem_dff.code_mem[1][4] ),
    .A2(_03355_),
    .B1(_03358_),
    .B2(\mem.mem_dff.code_mem[17][4] ),
    .C(_03356_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08271_ (.I(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08272_ (.A1(\mem.mem_dff.code_mem[5][4] ),
    .A2(_03352_),
    .B1(_03353_),
    .B2(\mem.mem_dff.code_mem[20][4] ),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08273_ (.A1(\mem.mem_dff.code_mem[2][4] ),
    .A2(_03349_),
    .B1(_03350_),
    .B2(\mem.mem_dff.code_mem[18][4] ),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08274_ (.A1(\mem.mem_dff.code_mem[19][4] ),
    .A2(_03366_),
    .B1(_03359_),
    .B2(\mem.mem_dff.code_mem[21][4] ),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08275_ (.A1(\mem.mem_dff.code_mem[3][4] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\mem.mem_dff.code_mem[4][4] ),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08276_ (.A1(_03464_),
    .A2(_03465_),
    .A3(_03466_),
    .A4(_03467_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08277_ (.A1(\mem.mem_dff.code_mem[16][4] ),
    .A2(_02536_),
    .B(_03463_),
    .C(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08278_ (.A1(\mem.mem_dff.code_mem[9][4] ),
    .A2(_03429_),
    .B1(_03430_),
    .B2(\mem.mem_dff.code_mem[28][4] ),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08279_ (.A1(\mem.mem_dff.code_mem[7][4] ),
    .A2(_03428_),
    .B1(_03432_),
    .B2(\mem.mem_dff.code_mem[14][4] ),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08280_ (.A1(_03461_),
    .A2(_03469_),
    .A3(_03470_),
    .A4(_03471_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08281_ (.I(_02015_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08282_ (.A1(\mem.mem_dff.code_mem[0][4] ),
    .A2(_03451_),
    .B1(_03456_),
    .B2(_03472_),
    .C(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08283_ (.I(_02986_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08284_ (.I(_02988_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08285_ (.A1(\mem.mem_dff.data_mem[2][4] ),
    .A2(_03043_),
    .B1(_03130_),
    .B2(\mem.mem_dff.data_mem[5][4] ),
    .C1(\mem.mem_dff.data_mem[7][4] ),
    .C2(_03321_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08286_ (.A1(\mem.mem_dff.data_mem[1][4] ),
    .A2(_03016_),
    .B1(_03070_),
    .B2(\mem.mem_dff.data_mem[3][4] ),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08287_ (.A1(\mem.mem_dff.data_mem[4][4] ),
    .A2(net227),
    .B1(_03329_),
    .B2(\mem.mem_dff.data_mem[6][4] ),
    .C(_03381_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08288_ (.A1(_03477_),
    .A2(_03478_),
    .A3(_03479_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08289_ (.A1(\mem.mem_dff.data_mem[0][4] ),
    .A2(_03475_),
    .B(_03476_),
    .C(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08290_ (.A1(_03474_),
    .A2(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08291_ (.I(_03335_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08292_ (.I0(\mem.dff_data_out[4] ),
    .I1(_03482_),
    .S(_03483_),
    .Z(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08293_ (.I(_03484_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08294_ (.A1(\mem.mem_dff.code_mem[15][5] ),
    .A2(_03368_),
    .B1(_03369_),
    .B2(\mem.mem_dff.code_mem[29][5] ),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08295_ (.A1(\mem.mem_dff.code_mem[6][5] ),
    .A2(_03388_),
    .B1(_03389_),
    .B2(\mem.mem_dff.code_mem[30][5] ),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08296_ (.A1(\mem.mem_dff.code_mem[23][5] ),
    .A2(_03391_),
    .B1(_03392_),
    .B2(\mem.mem_dff.code_mem[31][5] ),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08297_ (.A1(_03485_),
    .A2(_03486_),
    .A3(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08298_ (.A1(\mem.mem_dff.code_mem[8][5] ),
    .A2(_02293_),
    .B1(_02701_),
    .B2(\mem.mem_dff.code_mem[22][5] ),
    .C(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08299_ (.A1(\mem.mem_dff.code_mem[10][5] ),
    .A2(_03343_),
    .B1(_03344_),
    .B2(\mem.mem_dff.code_mem[24][5] ),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08300_ (.I(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08301_ (.A1(\mem.mem_dff.code_mem[25][5] ),
    .A2(_02789_),
    .B1(_02846_),
    .B2(\mem.mem_dff.code_mem[27][5] ),
    .C(_03491_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08302_ (.A1(\mem.mem_dff.code_mem[9][5] ),
    .A2(_03429_),
    .B1(_03432_),
    .B2(\mem.mem_dff.code_mem[14][5] ),
    .C1(\mem.mem_dff.code_mem[28][5] ),
    .C2(_03430_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08303_ (.A1(\mem.mem_dff.code_mem[7][5] ),
    .A2(_03428_),
    .B1(_02443_),
    .B2(\mem.mem_dff.code_mem[13][5] ),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08304_ (.A1(_03489_),
    .A2(_03492_),
    .A3(_03493_),
    .A4(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08305_ (.A1(\mem.mem_dff.code_mem[17][5] ),
    .A2(_02562_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08306_ (.A1(\mem.mem_dff.code_mem[1][5] ),
    .A2(_02071_),
    .B1(_03405_),
    .B2(\mem.mem_dff.code_mem[16][5] ),
    .C(_02027_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08307_ (.A1(\mem.mem_dff.code_mem[5][5] ),
    .A2(_03352_),
    .B1(_03353_),
    .B2(\mem.mem_dff.code_mem[20][5] ),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08308_ (.A1(\mem.mem_dff.code_mem[2][5] ),
    .A2(_03349_),
    .B1(_03350_),
    .B2(\mem.mem_dff.code_mem[18][5] ),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08309_ (.A1(\mem.mem_dff.code_mem[19][5] ),
    .A2(_03366_),
    .B1(_03359_),
    .B2(\mem.mem_dff.code_mem[21][5] ),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08310_ (.A1(\mem.mem_dff.code_mem[3][5] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\mem.mem_dff.code_mem[4][5] ),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08311_ (.A1(_03498_),
    .A2(_03499_),
    .A3(_03500_),
    .A4(_03501_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08312_ (.A1(\mem.mem_dff.code_mem[11][5] ),
    .A2(_03299_),
    .B1(_02414_),
    .B2(\mem.mem_dff.code_mem[12][5] ),
    .C1(\mem.mem_dff.code_mem[26][5] ),
    .C2(_03300_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08313_ (.A1(_03496_),
    .A2(_03497_),
    .A3(_03502_),
    .A4(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08314_ (.A1(\mem.mem_dff.code_mem[0][5] ),
    .A2(_03451_),
    .B1(_03495_),
    .B2(_03504_),
    .C(_03473_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08315_ (.A1(\mem.mem_dff.data_mem[1][5] ),
    .A2(_03016_),
    .B1(_03070_),
    .B2(\mem.mem_dff.data_mem[3][5] ),
    .C1(\mem.mem_dff.data_mem[7][5] ),
    .C2(_03321_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08316_ (.A1(\mem.mem_dff.data_mem[4][5] ),
    .A2(_03323_),
    .B1(_03324_),
    .B2(\mem.mem_dff.data_mem[5][5] ),
    .C(_03325_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08317_ (.A1(\mem.mem_dff.data_mem[2][5] ),
    .A2(_03327_),
    .B1(_03329_),
    .B2(\mem.mem_dff.data_mem[6][5] ),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08318_ (.A1(_03506_),
    .A2(_03507_),
    .A3(_03508_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08319_ (.A1(\mem.mem_dff.data_mem[0][5] ),
    .A2(_03475_),
    .B(_03476_),
    .C(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08320_ (.A1(_03505_),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08321_ (.I0(\mem.dff_data_out[5] ),
    .I1(_03511_),
    .S(_03483_),
    .Z(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08322_ (.I(_03512_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08323_ (.A1(\mem.mem_dff.code_mem[15][6] ),
    .A2(_03368_),
    .B1(_03369_),
    .B2(\mem.mem_dff.code_mem[29][6] ),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08324_ (.A1(\mem.mem_dff.code_mem[6][6] ),
    .A2(_03388_),
    .B1(_03389_),
    .B2(\mem.mem_dff.code_mem[30][6] ),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08325_ (.A1(\mem.mem_dff.code_mem[23][6] ),
    .A2(_03391_),
    .B1(_03392_),
    .B2(\mem.mem_dff.code_mem[31][6] ),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08326_ (.A1(_03513_),
    .A2(_03514_),
    .A3(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08327_ (.A1(\mem.mem_dff.code_mem[8][6] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\mem.mem_dff.code_mem[22][6] ),
    .C(_03516_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08328_ (.A1(\mem.mem_dff.code_mem[10][6] ),
    .A2(_03343_),
    .B1(_03344_),
    .B2(\mem.mem_dff.code_mem[24][6] ),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08329_ (.I(_03518_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08330_ (.A1(\mem.mem_dff.code_mem[25][6] ),
    .A2(_02789_),
    .B1(_02846_),
    .B2(\mem.mem_dff.code_mem[27][6] ),
    .C(_03519_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08331_ (.A1(\mem.mem_dff.code_mem[9][6] ),
    .A2(_02320_),
    .B1(_02468_),
    .B2(\mem.mem_dff.code_mem[14][6] ),
    .C1(\mem.mem_dff.code_mem[28][6] ),
    .C2(_03430_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08332_ (.A1(\mem.mem_dff.code_mem[7][6] ),
    .A2(_03428_),
    .B1(_02443_),
    .B2(\mem.mem_dff.code_mem[13][6] ),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08333_ (.A1(_03517_),
    .A2(_03520_),
    .A3(_03521_),
    .A4(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08334_ (.A1(\mem.mem_dff.code_mem[3][6] ),
    .A2(_02137_),
    .B1(_02173_),
    .B2(\mem.mem_dff.code_mem[4][6] ),
    .C1(\mem.mem_dff.code_mem[21][6] ),
    .C2(_02676_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08335_ (.A1(\mem.mem_dff.code_mem[5][6] ),
    .A2(_02200_),
    .B1(_02650_),
    .B2(\mem.mem_dff.code_mem[20][6] ),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08336_ (.A1(\mem.mem_dff.code_mem[2][6] ),
    .A2(_02098_),
    .B1(_02588_),
    .B2(\mem.mem_dff.code_mem[18][6] ),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08337_ (.A1(\mem.mem_dff.code_mem[1][6] ),
    .A2(_03355_),
    .B1(_03405_),
    .B2(\mem.mem_dff.code_mem[16][6] ),
    .C(_03356_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08338_ (.A1(\mem.mem_dff.code_mem[17][6] ),
    .A2(_03358_),
    .B1(_02620_),
    .B2(\mem.mem_dff.code_mem[19][6] ),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08339_ (.A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .A4(_03528_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _08340_ (.A1(\mem.mem_dff.code_mem[11][6] ),
    .A2(_03299_),
    .B1(_02415_),
    .B2(\mem.mem_dff.code_mem[12][6] ),
    .C1(\mem.mem_dff.code_mem[26][6] ),
    .C2(_03300_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08341_ (.A1(_03524_),
    .A2(_03529_),
    .A3(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08342_ (.A1(\mem.mem_dff.code_mem[0][6] ),
    .A2(_03451_),
    .B1(_03523_),
    .B2(_03531_),
    .C(_03473_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08343_ (.A1(\mem.mem_dff.data_mem[2][6] ),
    .A2(_03327_),
    .B1(_03375_),
    .B2(\mem.mem_dff.data_mem[6][6] ),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08344_ (.A1(\mem.mem_dff.data_mem[1][6] ),
    .A2(_03015_),
    .B1(_03069_),
    .B2(\mem.mem_dff.data_mem[3][6] ),
    .C1(\mem.mem_dff.data_mem[7][6] ),
    .C2(_03379_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08345_ (.A1(\mem.mem_dff.data_mem[4][6] ),
    .A2(_03323_),
    .B1(_03324_),
    .B2(\mem.mem_dff.data_mem[5][6] ),
    .C(_03325_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08346_ (.A1(_03533_),
    .A2(_03534_),
    .A3(_03535_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08347_ (.A1(\mem.mem_dff.data_mem[0][6] ),
    .A2(_03475_),
    .B(_03476_),
    .C(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08348_ (.A1(_03532_),
    .A2(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08349_ (.I0(\mem.dff_data_out[6] ),
    .I1(_03538_),
    .S(_03483_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08350_ (.I(_03539_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08351_ (.A1(\mem.mem_dff.code_mem[15][7] ),
    .A2(_02498_),
    .B1(_02901_),
    .B2(\mem.mem_dff.code_mem[29][7] ),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08352_ (.A1(\mem.mem_dff.code_mem[6][7] ),
    .A2(_02225_),
    .B1(_02926_),
    .B2(\mem.mem_dff.code_mem[30][7] ),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08353_ (.A1(\mem.mem_dff.code_mem[23][7] ),
    .A2(_02730_),
    .B1(_02956_),
    .B2(\mem.mem_dff.code_mem[31][7] ),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08354_ (.A1(_03540_),
    .A2(_03541_),
    .A3(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08355_ (.A1(\mem.mem_dff.code_mem[8][7] ),
    .A2(_03292_),
    .B1(_03293_),
    .B2(\mem.mem_dff.code_mem[22][7] ),
    .C(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08356_ (.A1(\mem.mem_dff.code_mem[10][7] ),
    .A2(_03343_),
    .B1(_03344_),
    .B2(\mem.mem_dff.code_mem[24][7] ),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08357_ (.I(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08358_ (.A1(\mem.mem_dff.code_mem[25][7] ),
    .A2(_03340_),
    .B1(_03341_),
    .B2(\mem.mem_dff.code_mem[27][7] ),
    .C(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08359_ (.A1(\mem.mem_dff.code_mem[7][7] ),
    .A2(_02257_),
    .B1(_03429_),
    .B2(\mem.mem_dff.code_mem[9][7] ),
    .C1(\mem.mem_dff.code_mem[28][7] ),
    .C2(_02875_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08360_ (.A1(\mem.mem_dff.code_mem[12][7] ),
    .A2(_02415_),
    .B1(_03432_),
    .B2(\mem.mem_dff.code_mem[14][7] ),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08361_ (.A1(_03544_),
    .A2(_03547_),
    .A3(_03548_),
    .A4(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08362_ (.A1(\mem.mem_dff.code_mem[16][7] ),
    .A2(_02536_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08363_ (.A1(\mem.mem_dff.code_mem[1][7] ),
    .A2(_02071_),
    .B1(_02562_),
    .B2(\mem.mem_dff.code_mem[17][7] ),
    .C(_02027_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08364_ (.A1(\mem.mem_dff.code_mem[5][7] ),
    .A2(_03352_),
    .B1(_03353_),
    .B2(\mem.mem_dff.code_mem[20][7] ),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08365_ (.A1(\mem.mem_dff.code_mem[2][7] ),
    .A2(_03349_),
    .B1(_03350_),
    .B2(\mem.mem_dff.code_mem[18][7] ),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08366_ (.A1(\mem.mem_dff.code_mem[19][7] ),
    .A2(_03366_),
    .B1(_03359_),
    .B2(\mem.mem_dff.code_mem[21][7] ),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08367_ (.A1(\mem.mem_dff.code_mem[3][7] ),
    .A2(_03364_),
    .B1(_03365_),
    .B2(\mem.mem_dff.code_mem[4][7] ),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08368_ (.A1(_03553_),
    .A2(_03554_),
    .A3(_03555_),
    .A4(_03556_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08369_ (.A1(\mem.mem_dff.code_mem[11][7] ),
    .A2(_02382_),
    .B1(_02442_),
    .B2(\mem.mem_dff.code_mem[13][7] ),
    .C1(\mem.mem_dff.code_mem[26][7] ),
    .C2(_02814_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08370_ (.A1(_03551_),
    .A2(_03552_),
    .A3(_03557_),
    .A4(_03558_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08371_ (.A1(\mem.mem_dff.code_mem[0][7] ),
    .A2(_03451_),
    .B1(_03550_),
    .B2(_03559_),
    .C(_03473_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08372_ (.A1(\mem.mem_dff.data_mem[1][7] ),
    .A2(_03377_),
    .B1(_03378_),
    .B2(\mem.mem_dff.data_mem[3][7] ),
    .C1(\mem.mem_dff.data_mem[7][7] ),
    .C2(_03321_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08373_ (.A1(\mem.mem_dff.data_mem[4][7] ),
    .A2(_03323_),
    .B1(_03324_),
    .B2(\mem.mem_dff.data_mem[5][7] ),
    .C(_03325_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08374_ (.A1(\mem.mem_dff.data_mem[2][7] ),
    .A2(_03327_),
    .B1(_03329_),
    .B2(\mem.mem_dff.data_mem[6][7] ),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08375_ (.A1(_03561_),
    .A2(_03562_),
    .A3(_03563_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08376_ (.A1(\mem.mem_dff.data_mem[0][7] ),
    .A2(_03475_),
    .B(_03476_),
    .C(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08377_ (.A1(_03560_),
    .A2(_03565_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08378_ (.I0(\mem.dff_data_out[7] ),
    .I1(_03566_),
    .S(_03483_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08379_ (.I(_03567_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08380_ (.I(_02003_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08381_ (.I(_03568_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08382_ (.A1(net253),
    .A2(_00763_),
    .A3(_01177_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08383_ (.A1(_02813_),
    .A2(_02986_),
    .A3(_03247_),
    .A4(_03570_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08384_ (.I(_03571_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08385_ (.I(_03572_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08386_ (.I(_03251_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08387_ (.A1(\mem.mem_io.past_write ),
    .A2(_03574_),
    .A3(_03570_),
    .B(_03571_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08388_ (.I(_03575_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08389_ (.A1(net120),
    .A2(_03573_),
    .B1(_03576_),
    .B2(_03073_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08390_ (.I(_03572_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08391_ (.I(_03575_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08392_ (.A1(net120),
    .A2(_02101_),
    .A3(_03578_),
    .A4(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08393_ (.A1(_03569_),
    .A2(_03577_),
    .A3(_03580_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08394_ (.I(_03568_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08395_ (.A1(net121),
    .A2(_03573_),
    .B1(_03576_),
    .B2(_03107_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08396_ (.A1(net121),
    .A2(_03107_),
    .A3(_03578_),
    .A4(_03579_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08397_ (.A1(_03581_),
    .A2(_03582_),
    .A3(_03583_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08398_ (.A1(net122),
    .A2(_03573_),
    .B1(_03576_),
    .B2(_03079_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08399_ (.A1(net122),
    .A2(_02108_),
    .A3(_03578_),
    .A4(_03579_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08400_ (.A1(_03581_),
    .A2(_03584_),
    .A3(_03585_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08401_ (.A1(net123),
    .A2(_03573_),
    .B1(_03576_),
    .B2(_03112_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08402_ (.A1(net123),
    .A2(_03112_),
    .A3(_03578_),
    .A4(_03579_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08403_ (.A1(_03581_),
    .A2(_03586_),
    .A3(_03587_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08404_ (.I(_03572_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08405_ (.I(_03575_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08406_ (.A1(net124),
    .A2(_03588_),
    .B1(_03589_),
    .B2(_03086_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08407_ (.I(_03572_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08408_ (.I(_03575_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08409_ (.A1(net124),
    .A2(_02116_),
    .A3(_03591_),
    .A4(_03592_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08410_ (.A1(_03581_),
    .A2(_03590_),
    .A3(_03593_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08411_ (.I(_03568_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08412_ (.A1(net125),
    .A2(_03588_),
    .B1(_03589_),
    .B2(_03090_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08413_ (.A1(net125),
    .A2(_02121_),
    .A3(_03591_),
    .A4(_03592_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08414_ (.A1(_03594_),
    .A2(_03595_),
    .A3(_03596_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08415_ (.A1(net126),
    .A2(_03588_),
    .B1(_03589_),
    .B2(_03122_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08416_ (.A1(net126),
    .A2(_03122_),
    .A3(_03591_),
    .A4(_03592_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08417_ (.A1(_03594_),
    .A2(_03597_),
    .A3(_03598_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08418_ (.A1(net127),
    .A2(_03588_),
    .B1(_03589_),
    .B2(_03125_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08419_ (.A1(net127),
    .A2(_03125_),
    .A3(_03591_),
    .A4(_03592_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08420_ (.A1(_03594_),
    .A2(_03599_),
    .A3(_03600_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08421_ (.A1(_02985_),
    .A2(_02256_),
    .A3(_03248_),
    .A4(_03570_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08422_ (.I(_03601_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08423_ (.I(_03601_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08424_ (.A1(net112),
    .A2(_03603_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08425_ (.I(_02009_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08426_ (.A1(_02031_),
    .A2(_03602_),
    .B(_03604_),
    .C(_03605_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08427_ (.A1(net113),
    .A2(_03603_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08428_ (.A1(_02037_),
    .A2(_03602_),
    .B(_03606_),
    .C(_03605_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08429_ (.A1(net114),
    .A2(_03603_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08430_ (.A1(_02041_),
    .A2(_03602_),
    .B(_03607_),
    .C(_03605_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(net115),
    .A2(_03603_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08432_ (.A1(_02045_),
    .A2(_03602_),
    .B(_03608_),
    .C(_03605_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08433_ (.I(_03601_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08434_ (.I(_03601_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08435_ (.A1(net116),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08436_ (.I(_02009_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08437_ (.A1(_02051_),
    .A2(_03609_),
    .B(_03611_),
    .C(_03612_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08438_ (.A1(net117),
    .A2(_03610_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08439_ (.A1(_02056_),
    .A2(_03609_),
    .B(_03613_),
    .C(_03612_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08440_ (.A1(net118),
    .A2(_03610_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08441_ (.A1(_02060_),
    .A2(_03609_),
    .B(_03614_),
    .C(_03612_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08442_ (.A1(net119),
    .A2(_03610_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08443_ (.A1(_02064_),
    .A2(_03609_),
    .B(_03615_),
    .C(_03612_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08444_ (.A1(_03282_),
    .A2(_03244_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08445_ (.I(_01660_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08446_ (.A1(_01662_),
    .A2(_01663_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(_01664_),
    .A2(_03617_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08448_ (.A1(_03616_),
    .A2(_01696_),
    .A3(_03618_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08449_ (.I(_01630_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08450_ (.I(_03620_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08451_ (.I(_03621_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08452_ (.I(_01769_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08453_ (.A1(_03622_),
    .A2(_03623_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08454_ (.I(_01631_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08455_ (.A1(_03625_),
    .A2(_01243_),
    .B(\intr[1] ),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08456_ (.I(_03568_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08457_ (.A1(_03619_),
    .A2(_03624_),
    .B(_03626_),
    .C(_03627_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08458_ (.I(_01604_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08459_ (.I(_01588_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08460_ (.A1(_03629_),
    .A2(_03194_),
    .A3(_03195_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08461_ (.A1(_03628_),
    .A2(_03199_),
    .A3(_01637_),
    .A4(_03630_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08462_ (.I(_03631_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08463_ (.I(_01757_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08464_ (.I0(_01673_),
    .I1(_01651_),
    .S(_01679_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08465_ (.I(_03634_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08466_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08467_ (.I(_01684_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08468_ (.A1(_01689_),
    .A2(_01693_),
    .A3(_01698_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08469_ (.A1(_03638_),
    .A2(_01703_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08470_ (.A1(_01711_),
    .A2(_03639_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08471_ (.A1(_03636_),
    .A2(_03637_),
    .A3(_01692_),
    .A4(_03640_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08472_ (.I(_03641_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08473_ (.A1(_03629_),
    .A2(_03194_),
    .A3(_03195_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08474_ (.A1(_03628_),
    .A2(_03199_),
    .A3(_01636_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08475_ (.I(_03644_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08476_ (.A1(_03643_),
    .A2(_03645_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08477_ (.A1(_03185_),
    .A2(_03641_),
    .A3(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08478_ (.I(_03647_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08479_ (.A1(_03633_),
    .A2(_03642_),
    .B1(_03648_),
    .B2(\stack[19][0] ),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08480_ (.A1(_01183_),
    .A2(_03632_),
    .B(_03649_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08481_ (.I(_03214_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08482_ (.A1(_03650_),
    .A2(_03642_),
    .B1(_03648_),
    .B2(\stack[19][1] ),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08483_ (.A1(_01764_),
    .A2(_03632_),
    .B(_03651_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08484_ (.I(_03217_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08485_ (.A1(_03652_),
    .A2(_03642_),
    .B1(_03648_),
    .B2(\stack[19][2] ),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08486_ (.A1(_01797_),
    .A2(_03632_),
    .B(_03653_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08487_ (.I(_03220_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08488_ (.A1(_03654_),
    .A2(_03642_),
    .B1(_03648_),
    .B2(\stack[19][3] ),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08489_ (.A1(_01829_),
    .A2(_03632_),
    .B(_03655_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08490_ (.I(_03223_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08491_ (.I(_03647_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08492_ (.A1(_03656_),
    .A2(_03641_),
    .B1(_03657_),
    .B2(\stack[19][4] ),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08493_ (.A1(_01861_),
    .A2(_03631_),
    .B(_03658_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08494_ (.I(_03227_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08495_ (.A1(_03659_),
    .A2(_03641_),
    .B1(_03657_),
    .B2(\stack[19][5] ),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08496_ (.A1(_01893_),
    .A2(_03631_),
    .B(_03660_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_03636_),
    .A2(_01925_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08498_ (.A1(_01931_),
    .A2(_03661_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08499_ (.I(_03640_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08500_ (.I(_03663_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08501_ (.A1(_03662_),
    .A2(_03664_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08502_ (.A1(_03238_),
    .A2(_03646_),
    .B1(_03657_),
    .B2(\stack[19][6] ),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08503_ (.A1(_01964_),
    .A2(_03665_),
    .B(_03666_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08504_ (.A1(net152),
    .A2(_03646_),
    .B1(_03657_),
    .B2(\stack[19][7] ),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08505_ (.A1(_01991_),
    .A2(_03665_),
    .B(_03667_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08506_ (.A1(_03628_),
    .A2(_01707_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08507_ (.A1(_03668_),
    .A2(_01637_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08508_ (.A1(_03198_),
    .A2(_03669_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08509_ (.I(_03670_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08510_ (.I(_01675_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08511_ (.I(_03187_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08512_ (.A1(_03638_),
    .A2(_01703_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08513_ (.A1(_03191_),
    .A2(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08514_ (.A1(_03672_),
    .A2(_03673_),
    .A3(_03189_),
    .A4(_03675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08515_ (.I(_03676_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08516_ (.A1(_01707_),
    .A2(_03200_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08517_ (.I(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08518_ (.A1(_03198_),
    .A2(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08519_ (.A1(_03185_),
    .A2(_03676_),
    .A3(_03680_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08520_ (.I(_03681_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08521_ (.A1(_03633_),
    .A2(_03677_),
    .B1(_03682_),
    .B2(\stack[29][0] ),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08522_ (.A1(_01183_),
    .A2(_03671_),
    .B(_03683_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08523_ (.A1(_03650_),
    .A2(_03677_),
    .B1(_03682_),
    .B2(\stack[29][1] ),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08524_ (.A1(_01764_),
    .A2(_03671_),
    .B(_03684_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08525_ (.A1(_03652_),
    .A2(_03677_),
    .B1(_03682_),
    .B2(\stack[29][2] ),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08526_ (.A1(_01797_),
    .A2(_03671_),
    .B(_03685_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08527_ (.A1(_03654_),
    .A2(_03677_),
    .B1(_03682_),
    .B2(\stack[29][3] ),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08528_ (.A1(_01829_),
    .A2(_03671_),
    .B(_03686_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08529_ (.I(_03681_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08530_ (.A1(_03656_),
    .A2(_03676_),
    .B1(_03687_),
    .B2(\stack[29][4] ),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08531_ (.A1(_01861_),
    .A2(_03670_),
    .B(_03688_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08532_ (.A1(_03659_),
    .A2(_03676_),
    .B1(_03687_),
    .B2(\stack[29][5] ),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08533_ (.A1(_01893_),
    .A2(_03670_),
    .B(_03689_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08534_ (.A1(_01711_),
    .A2(_03674_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08535_ (.I(_03690_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08536_ (.I(_03691_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08537_ (.A1(_03232_),
    .A2(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08538_ (.I(_03237_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08539_ (.A1(_03694_),
    .A2(_03680_),
    .B1(_03687_),
    .B2(\stack[29][6] ),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08540_ (.A1(_01964_),
    .A2(_03693_),
    .B(_03695_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08541_ (.I(_01170_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08542_ (.A1(_03696_),
    .A2(_03680_),
    .B1(_03687_),
    .B2(\stack[29][7] ),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08543_ (.A1(_01991_),
    .A2(_03693_),
    .B(_03697_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08544_ (.I(_03645_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08545_ (.A1(_03194_),
    .A2(_03195_),
    .A3(_03197_),
    .A4(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08546_ (.I(_03699_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08547_ (.I(_01683_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08548_ (.A1(_03191_),
    .A2(_03639_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08549_ (.A1(_01676_),
    .A2(_03701_),
    .A3(_01691_),
    .A4(_03702_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08550_ (.I(_03703_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08551_ (.A1(_03167_),
    .A2(_03704_),
    .A3(_03699_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08552_ (.I(_03705_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08553_ (.I(_03703_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_03633_),
    .A2(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08555_ (.A1(_01182_),
    .A2(_03700_),
    .B1(_03706_),
    .B2(_01326_),
    .C(_03708_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08556_ (.I(\stack[31][1] ),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08557_ (.A1(_03215_),
    .A2(_03707_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08558_ (.A1(_01763_),
    .A2(_03700_),
    .B1(_03705_),
    .B2(_03709_),
    .C(_03710_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08559_ (.I(_03707_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08560_ (.I(_01795_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08561_ (.A1(_03712_),
    .A2(_03700_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08562_ (.A1(_03218_),
    .A2(_03711_),
    .B(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08563_ (.A1(_01315_),
    .A2(_03706_),
    .B(_03714_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08564_ (.I(\stack[31][3] ),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08565_ (.I(_01827_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08566_ (.I(_03699_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08567_ (.A1(_03716_),
    .A2(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08568_ (.A1(_03221_),
    .A2(_03711_),
    .B(_03718_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08569_ (.A1(_03715_),
    .A2(_03706_),
    .B(_03719_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08570_ (.I(\stack[31][4] ),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08571_ (.I(_01859_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08572_ (.A1(_03721_),
    .A2(_03717_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08573_ (.A1(_03224_),
    .A2(_03711_),
    .B(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08574_ (.A1(_03720_),
    .A2(_03706_),
    .B(_03723_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08575_ (.I(_03227_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08576_ (.A1(_03724_),
    .A2(_03711_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08577_ (.A1(_01999_),
    .A2(_03699_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08578_ (.A1(_03707_),
    .A2(_03726_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08579_ (.I(_01891_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08580_ (.A1(_03728_),
    .A2(_03700_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08581_ (.A1(\stack[31][5] ),
    .A2(_03727_),
    .B(_03729_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_03725_),
    .A2(_03730_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08583_ (.I(_01962_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08584_ (.I(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_01937_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08586_ (.A1(_03733_),
    .A2(_03717_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08587_ (.A1(\stack[31][6] ),
    .A2(_03727_),
    .B(_03734_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08588_ (.A1(_03732_),
    .A2(_03704_),
    .B(_03735_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08589_ (.I(_01990_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08590_ (.I(_01975_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08591_ (.A1(_03737_),
    .A2(_03717_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08592_ (.A1(\stack[31][7] ),
    .A2(_03727_),
    .B(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08593_ (.A1(_03736_),
    .A2(_03704_),
    .B(_03739_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08594_ (.I(_02002_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08595_ (.I(_01676_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08596_ (.A1(_03741_),
    .A2(_01685_),
    .A3(_01692_),
    .A4(_03640_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08597_ (.I(_03644_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08598_ (.A1(_01618_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08599_ (.A1(_03740_),
    .A2(_03742_),
    .A3(_03744_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08600_ (.I(_03745_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08601_ (.A1(\stack[3][0] ),
    .A2(_03746_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08602_ (.I(_03742_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08603_ (.I(_03744_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08604_ (.A1(_03208_),
    .A2(_03748_),
    .B1(_03749_),
    .B2(net144),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(_03747_),
    .A2(_03750_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08606_ (.A1(\stack[3][1] ),
    .A2(_03746_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08607_ (.I(_03214_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08608_ (.A1(_03752_),
    .A2(_03748_),
    .B1(_03749_),
    .B2(net145),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08609_ (.A1(_03751_),
    .A2(_03753_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(\stack[3][2] ),
    .A2(_03746_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08611_ (.I(_03217_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08612_ (.A1(_03755_),
    .A2(_03748_),
    .B1(_03749_),
    .B2(net146),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08613_ (.A1(_03754_),
    .A2(_03756_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08614_ (.A1(\stack[3][3] ),
    .A2(_03746_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08615_ (.I(_03220_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08616_ (.A1(_03758_),
    .A2(_03742_),
    .B1(_03749_),
    .B2(net147),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08617_ (.A1(_03757_),
    .A2(_03759_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08618_ (.I(_03745_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08619_ (.A1(\stack[3][4] ),
    .A2(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08620_ (.I(_03223_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08621_ (.I(_03744_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08622_ (.A1(_03762_),
    .A2(_03742_),
    .B1(_03763_),
    .B2(net148),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08623_ (.A1(_03761_),
    .A2(_03764_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08624_ (.A1(_03724_),
    .A2(_03748_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08625_ (.A1(net149),
    .A2(_03763_),
    .B1(_03760_),
    .B2(\stack[3][5] ),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08626_ (.A1(_03765_),
    .A2(_03766_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08627_ (.A1(_01932_),
    .A2(_03664_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08628_ (.A1(_03694_),
    .A2(_03763_),
    .B1(_03760_),
    .B2(\stack[3][6] ),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08629_ (.A1(_03732_),
    .A2(_03767_),
    .B(_03768_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08630_ (.A1(_03696_),
    .A2(_03763_),
    .B1(_03760_),
    .B2(\stack[3][7] ),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08631_ (.A1(_03736_),
    .A2(_03767_),
    .B(_03769_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08632_ (.A1(_01598_),
    .A2(_01604_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08633_ (.I(_01616_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08634_ (.A1(_01588_),
    .A2(_03770_),
    .A3(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08635_ (.A1(_03201_),
    .A2(_03772_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08636_ (.I(_03773_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(_03774_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08638_ (.I(_01757_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(_01929_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08640_ (.A1(_03741_),
    .A2(_03637_),
    .A3(_03777_),
    .A4(_03234_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08641_ (.I(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08642_ (.I(_01643_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(_03780_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08644_ (.A1(_03781_),
    .A2(_03778_),
    .A3(_03773_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08645_ (.I(_03782_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08646_ (.A1(_03776_),
    .A2(_03779_),
    .B1(_03783_),
    .B2(\stack[4][0] ),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08647_ (.A1(_01183_),
    .A2(_03775_),
    .B(_03784_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08648_ (.I(_01763_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08649_ (.A1(_03650_),
    .A2(_03779_),
    .B1(_03783_),
    .B2(\stack[4][1] ),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08650_ (.A1(_03785_),
    .A2(_03775_),
    .B(_03786_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08651_ (.I(_01796_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08652_ (.A1(_03652_),
    .A2(_03779_),
    .B1(_03783_),
    .B2(\stack[4][2] ),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08653_ (.A1(_03787_),
    .A2(_03775_),
    .B(_03788_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08654_ (.I(_01828_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08655_ (.A1(_03654_),
    .A2(_03779_),
    .B1(_03783_),
    .B2(\stack[4][3] ),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08656_ (.A1(_03789_),
    .A2(_03775_),
    .B(_03790_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08657_ (.I(_01860_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08658_ (.I(_03782_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08659_ (.A1(_03656_),
    .A2(_03778_),
    .B1(_03792_),
    .B2(\stack[4][4] ),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08660_ (.A1(_03791_),
    .A2(_03774_),
    .B(_03793_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08661_ (.I(_01892_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08662_ (.A1(_03659_),
    .A2(_03778_),
    .B1(_03792_),
    .B2(\stack[4][5] ),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08663_ (.A1(_03794_),
    .A2(_03774_),
    .B(_03795_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08664_ (.A1(_01926_),
    .A2(_03230_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(_03235_),
    .A2(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08666_ (.A1(_03694_),
    .A2(_03773_),
    .B1(_03792_),
    .B2(\stack[4][6] ),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08667_ (.A1(_03732_),
    .A2(_03797_),
    .B(_03798_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08668_ (.A1(_03696_),
    .A2(_03773_),
    .B1(_03792_),
    .B2(\stack[4][7] ),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08669_ (.A1(_03736_),
    .A2(_03797_),
    .B(_03799_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08670_ (.A1(_03741_),
    .A2(_03637_),
    .A3(_03777_),
    .A4(_03691_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08671_ (.A1(_03679_),
    .A2(_03772_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08672_ (.A1(_03781_),
    .A2(_03800_),
    .A3(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08673_ (.I(_03802_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08674_ (.A1(\stack[5][0] ),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08675_ (.I(_03800_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08676_ (.A1(_03208_),
    .A2(_03805_),
    .B1(_03801_),
    .B2(net144),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08677_ (.A1(_03804_),
    .A2(_03806_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08678_ (.I(_03772_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08679_ (.A1(_03669_),
    .A2(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08680_ (.I(_03808_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08681_ (.A1(_03650_),
    .A2(_03805_),
    .B1(_03803_),
    .B2(\stack[5][1] ),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08682_ (.A1(_03785_),
    .A2(_03809_),
    .B(_03810_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08683_ (.A1(_03652_),
    .A2(_03805_),
    .B1(_03803_),
    .B2(\stack[5][2] ),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08684_ (.A1(_03787_),
    .A2(_03809_),
    .B(_03811_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08685_ (.A1(_03654_),
    .A2(_03805_),
    .B1(_03803_),
    .B2(\stack[5][3] ),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08686_ (.A1(_03789_),
    .A2(_03809_),
    .B(_03812_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08687_ (.I(_03802_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08688_ (.A1(_03656_),
    .A2(_03800_),
    .B1(_03813_),
    .B2(\stack[5][4] ),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03791_),
    .A2(_03809_),
    .B(_03814_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08690_ (.A1(_03659_),
    .A2(_03800_),
    .B1(_03813_),
    .B2(\stack[5][5] ),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08691_ (.A1(_03794_),
    .A2(_03808_),
    .B(_03815_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08692_ (.A1(_03692_),
    .A2(_03796_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08693_ (.A1(_03694_),
    .A2(_03801_),
    .B1(_03813_),
    .B2(\stack[5][6] ),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08694_ (.A1(_03732_),
    .A2(_03816_),
    .B(_03817_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08695_ (.A1(_03696_),
    .A2(_03801_),
    .B1(_03813_),
    .B2(\stack[5][7] ),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08696_ (.A1(_03736_),
    .A2(_03816_),
    .B(_03818_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08697_ (.I(_01182_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08698_ (.I(_03201_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08699_ (.A1(_01587_),
    .A2(_03196_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08700_ (.A1(_03770_),
    .A2(_03771_),
    .A3(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08701_ (.I(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08702_ (.I(_03823_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08703_ (.A1(_03820_),
    .A2(_03824_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08704_ (.I(_03825_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08705_ (.I(_03634_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08706_ (.I(_01929_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08707_ (.A1(_03827_),
    .A2(_03673_),
    .A3(_03828_),
    .A4(_03192_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08708_ (.I(_03829_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08709_ (.A1(_03820_),
    .A2(_03823_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08710_ (.A1(_03781_),
    .A2(_03829_),
    .A3(_03831_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08711_ (.I(_03832_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08712_ (.A1(_03776_),
    .A2(_03830_),
    .B1(_03833_),
    .B2(\stack[8][0] ),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08713_ (.A1(_03819_),
    .A2(_03826_),
    .B(_03834_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08714_ (.I(_03214_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08715_ (.A1(_03835_),
    .A2(_03830_),
    .B1(_03833_),
    .B2(\stack[8][1] ),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08716_ (.A1(_03785_),
    .A2(_03826_),
    .B(_03836_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08717_ (.I(_03217_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08718_ (.A1(_03837_),
    .A2(_03830_),
    .B1(_03833_),
    .B2(\stack[8][2] ),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08719_ (.A1(_03787_),
    .A2(_03826_),
    .B(_03838_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08720_ (.I(_03220_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08721_ (.I(_03832_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08722_ (.A1(_03839_),
    .A2(_03830_),
    .B1(_03840_),
    .B2(\stack[8][3] ),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08723_ (.A1(_03789_),
    .A2(_03826_),
    .B(_03841_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08724_ (.I(_03223_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08725_ (.A1(_03842_),
    .A2(_03829_),
    .B1(_03840_),
    .B2(\stack[8][4] ),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08726_ (.A1(_03791_),
    .A2(_03825_),
    .B(_03843_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08727_ (.I(_03227_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08728_ (.A1(_03844_),
    .A2(_03829_),
    .B1(_03840_),
    .B2(\stack[8][5] ),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08729_ (.A1(_03794_),
    .A2(_03825_),
    .B(_03845_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08730_ (.I(_03731_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08731_ (.I(_03234_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08732_ (.A1(_03636_),
    .A2(_01925_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08733_ (.A1(_01931_),
    .A2(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(_03847_),
    .A2(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08735_ (.I(_03237_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08736_ (.A1(_03851_),
    .A2(_03831_),
    .B1(_03840_),
    .B2(\stack[8][6] ),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08737_ (.A1(_03846_),
    .A2(_03850_),
    .B(_03852_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08738_ (.I(_01989_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08739_ (.I(_03853_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08740_ (.I(_03737_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08741_ (.I(_03855_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08742_ (.A1(\stack[8][7] ),
    .A2(_03833_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08743_ (.A1(_03854_),
    .A2(_03850_),
    .B1(_03825_),
    .B2(_03856_),
    .C(_03857_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08744_ (.I(_03634_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08745_ (.A1(_03858_),
    .A2(_03188_),
    .A3(_03828_),
    .A4(_03702_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08746_ (.A1(_03743_),
    .A2(_03823_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08747_ (.A1(_03740_),
    .A2(_03859_),
    .A3(_03860_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08748_ (.I(_03861_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(\stack[11][0] ),
    .A2(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08750_ (.I(_03859_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08751_ (.I(_03860_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08752_ (.I(_00842_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08753_ (.A1(_03208_),
    .A2(_03864_),
    .B1(_03865_),
    .B2(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08754_ (.A1(_03863_),
    .A2(_03867_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08755_ (.I(_01762_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08756_ (.I(_03868_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08757_ (.I(_03645_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08758_ (.A1(_03870_),
    .A2(_03824_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08759_ (.I(_03861_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08760_ (.A1(\stack[11][1] ),
    .A2(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_03752_),
    .A2(_03864_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08762_ (.A1(_03869_),
    .A2(_03871_),
    .B(_03873_),
    .C(_03874_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08763_ (.A1(\stack[11][2] ),
    .A2(_03862_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08764_ (.A1(_03755_),
    .A2(_03864_),
    .B1(_03865_),
    .B2(net146),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(_03875_),
    .A2(_03876_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08766_ (.A1(\stack[11][3] ),
    .A2(_03862_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08767_ (.A1(_03758_),
    .A2(_03859_),
    .B1(_03865_),
    .B2(net147),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(_03877_),
    .A2(_03878_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08769_ (.I(_03721_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08770_ (.A1(\stack[11][4] ),
    .A2(_03872_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08771_ (.A1(_03762_),
    .A2(_03864_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08772_ (.A1(_03879_),
    .A2(_03871_),
    .B(_03880_),
    .C(_03881_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08773_ (.I(_03728_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08774_ (.A1(_03228_),
    .A2(_03859_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08775_ (.A1(\stack[11][5] ),
    .A2(_03862_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08776_ (.A1(_03882_),
    .A2(_03871_),
    .B(_03883_),
    .C(_03884_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08777_ (.A1(_03664_),
    .A2(_03849_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08778_ (.A1(_03851_),
    .A2(_03865_),
    .B1(_03872_),
    .B2(\stack[11][6] ),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_03846_),
    .A2(_03885_),
    .B(_03886_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08780_ (.I(_03853_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(\stack[11][7] ),
    .A2(_03872_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08782_ (.A1(_03887_),
    .A2(_03885_),
    .B1(_03871_),
    .B2(_03856_),
    .C(_03888_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08783_ (.I(_01181_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08784_ (.I(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08785_ (.A1(_01639_),
    .A2(_03807_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08786_ (.I(_03891_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08787_ (.A1(_01677_),
    .A2(_01685_),
    .A3(_01930_),
    .A4(_01713_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08788_ (.A1(_01639_),
    .A2(_03807_),
    .B(_02008_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08789_ (.A1(_03893_),
    .A2(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08790_ (.I(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(\stack[6][0] ),
    .A2(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08792_ (.I(_03207_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08793_ (.I(_03893_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08794_ (.A1(_03898_),
    .A2(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08795_ (.A1(_03890_),
    .A2(_03892_),
    .B(_03897_),
    .C(_03900_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08796_ (.I(_03891_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08797_ (.A1(_03835_),
    .A2(_03899_),
    .B1(_03896_),
    .B2(\stack[6][1] ),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08798_ (.A1(_03785_),
    .A2(_03901_),
    .B(_03902_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08799_ (.I(_03895_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08800_ (.A1(_03837_),
    .A2(_03899_),
    .B1(_03903_),
    .B2(\stack[6][2] ),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08801_ (.A1(_03787_),
    .A2(_03901_),
    .B(_03904_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(_03839_),
    .A2(_03899_),
    .B1(_03903_),
    .B2(\stack[6][3] ),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08803_ (.A1(_03789_),
    .A2(_03901_),
    .B(_03905_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08804_ (.A1(_03842_),
    .A2(_03893_),
    .B1(_03903_),
    .B2(\stack[6][4] ),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08805_ (.A1(_03791_),
    .A2(_03901_),
    .B(_03906_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08806_ (.A1(_03844_),
    .A2(_03893_),
    .B1(_03903_),
    .B2(\stack[6][5] ),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08807_ (.A1(_03794_),
    .A2(_03892_),
    .B(_03907_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08808_ (.I(_01963_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08809_ (.I(_01713_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08810_ (.A1(_03909_),
    .A2(_03796_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08811_ (.A1(\stack[6][6] ),
    .A2(_03896_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08812_ (.A1(_03908_),
    .A2(_03910_),
    .B1(_03892_),
    .B2(_03733_),
    .C(_03911_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08813_ (.A1(\stack[6][7] ),
    .A2(_03896_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08814_ (.A1(_03887_),
    .A2(_03910_),
    .B1(_03892_),
    .B2(_03856_),
    .C(_03912_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08815_ (.A1(_03741_),
    .A2(_03637_),
    .A3(_01930_),
    .A4(_03640_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08816_ (.A1(_03645_),
    .A2(_03807_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08817_ (.A1(_03185_),
    .A2(_03913_),
    .A3(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08818_ (.I(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08819_ (.A1(\stack[7][0] ),
    .A2(_03916_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08820_ (.I(_03207_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08821_ (.I(_03913_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08822_ (.I(_03914_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08823_ (.A1(_03918_),
    .A2(_03919_),
    .B1(_03920_),
    .B2(_03866_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(_03917_),
    .A2(_03921_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08825_ (.A1(\stack[7][1] ),
    .A2(_03916_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08826_ (.A1(_03215_),
    .A2(_03919_),
    .B1(_03920_),
    .B2(net145),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(_03922_),
    .A2(_03923_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08828_ (.A1(\stack[7][2] ),
    .A2(_03916_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08829_ (.A1(_03755_),
    .A2(_03919_),
    .B1(_03920_),
    .B2(net146),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08830_ (.A1(_03924_),
    .A2(_03925_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08831_ (.A1(\stack[7][3] ),
    .A2(_03916_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08832_ (.A1(_03758_),
    .A2(_03913_),
    .B1(_03920_),
    .B2(net147),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(_03926_),
    .A2(_03927_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08834_ (.I(_03915_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(\stack[7][4] ),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08836_ (.I(_03914_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08837_ (.A1(_03224_),
    .A2(_03913_),
    .B1(_03930_),
    .B2(net148),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08838_ (.A1(_03929_),
    .A2(_03931_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(_03724_),
    .A2(_03919_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08840_ (.A1(net149),
    .A2(_03930_),
    .B1(_03928_),
    .B2(\stack[7][5] ),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08841_ (.A1(_03932_),
    .A2(_03933_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08842_ (.A1(_03664_),
    .A2(_03796_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08843_ (.A1(_03851_),
    .A2(_03930_),
    .B1(_03928_),
    .B2(\stack[7][6] ),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08844_ (.A1(_03846_),
    .A2(_03934_),
    .B(_03935_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08845_ (.I(_01990_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08846_ (.I(_01170_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08847_ (.A1(_03937_),
    .A2(_03930_),
    .B1(_03928_),
    .B2(\stack[7][7] ),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08848_ (.A1(_03936_),
    .A2(_03934_),
    .B(_03938_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08849_ (.A1(_03770_),
    .A2(_03771_),
    .A3(_03197_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08850_ (.I(_03939_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08851_ (.I(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08852_ (.A1(_01640_),
    .A2(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08853_ (.I(_03942_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08854_ (.I(_01928_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08855_ (.A1(_01704_),
    .A2(_03191_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08856_ (.A1(_03672_),
    .A2(_03673_),
    .A3(_03944_),
    .A4(_03945_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08857_ (.I(_03946_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08858_ (.A1(_01639_),
    .A2(_03940_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08859_ (.A1(_03781_),
    .A2(_03946_),
    .A3(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08860_ (.I(_03949_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08861_ (.A1(_03776_),
    .A2(_03947_),
    .B1(_03950_),
    .B2(\stack[26][0] ),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08862_ (.A1(_03819_),
    .A2(_03943_),
    .B(_03951_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08863_ (.I(_01763_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08864_ (.A1(_03835_),
    .A2(_03947_),
    .B1(_03950_),
    .B2(\stack[26][1] ),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08865_ (.A1(_03952_),
    .A2(_03943_),
    .B(_03953_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08866_ (.I(_01796_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08867_ (.I(_03949_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08868_ (.A1(_03837_),
    .A2(_03947_),
    .B1(_03955_),
    .B2(\stack[26][2] ),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08869_ (.A1(_03954_),
    .A2(_03943_),
    .B(_03956_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08870_ (.I(_01828_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08871_ (.A1(_03839_),
    .A2(_03947_),
    .B1(_03955_),
    .B2(\stack[26][3] ),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08872_ (.A1(_03957_),
    .A2(_03943_),
    .B(_03958_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08873_ (.I(_01860_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08874_ (.A1(_03842_),
    .A2(_03946_),
    .B1(_03955_),
    .B2(\stack[26][4] ),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08875_ (.A1(_03959_),
    .A2(_03942_),
    .B(_03960_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08876_ (.I(_01892_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08877_ (.A1(_03844_),
    .A2(_03946_),
    .B1(_03955_),
    .B2(\stack[26][5] ),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08878_ (.A1(_03961_),
    .A2(_03942_),
    .B(_03962_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08879_ (.I(_01963_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08880_ (.A1(_01931_),
    .A2(_03231_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(_01933_),
    .A2(_03964_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08882_ (.A1(\stack[26][6] ),
    .A2(_03950_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08883_ (.A1(net151),
    .A2(_03948_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08884_ (.A1(_03963_),
    .A2(_03965_),
    .B(_03966_),
    .C(_03967_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(\stack[26][7] ),
    .A2(_03950_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08886_ (.A1(_03887_),
    .A2(_03965_),
    .B1(_03942_),
    .B2(_03856_),
    .C(_03968_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08887_ (.A1(_01640_),
    .A2(_03824_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08888_ (.I(_03969_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08889_ (.A1(_03827_),
    .A2(_03673_),
    .A3(_03944_),
    .A4(_03945_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08890_ (.I(_03971_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08891_ (.I(_03780_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08892_ (.A1(_01715_),
    .A2(_03823_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08893_ (.A1(_03973_),
    .A2(_03971_),
    .A3(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08894_ (.I(_03975_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08895_ (.A1(_03776_),
    .A2(_03972_),
    .B1(_03976_),
    .B2(\stack[10][0] ),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08896_ (.A1(_03819_),
    .A2(_03970_),
    .B(_03977_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08897_ (.A1(_03835_),
    .A2(_03972_),
    .B1(_03976_),
    .B2(\stack[10][1] ),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08898_ (.A1(_03952_),
    .A2(_03970_),
    .B(_03978_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08899_ (.I(_03975_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08900_ (.A1(_03837_),
    .A2(_03972_),
    .B1(_03979_),
    .B2(\stack[10][2] ),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08901_ (.A1(_03954_),
    .A2(_03970_),
    .B(_03980_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08902_ (.A1(_03839_),
    .A2(_03972_),
    .B1(_03979_),
    .B2(\stack[10][3] ),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08903_ (.A1(_03957_),
    .A2(_03970_),
    .B(_03981_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08904_ (.A1(_03842_),
    .A2(_03971_),
    .B1(_03979_),
    .B2(\stack[10][4] ),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08905_ (.A1(_03959_),
    .A2(_03969_),
    .B(_03982_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08906_ (.A1(_03844_),
    .A2(_03971_),
    .B1(_03979_),
    .B2(\stack[10][5] ),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08907_ (.A1(_03961_),
    .A2(_03969_),
    .B(_03983_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(_01933_),
    .A2(_03849_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(\stack[10][6] ),
    .A2(_03976_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(net151),
    .A2(_03974_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08911_ (.A1(_03963_),
    .A2(_03984_),
    .B(_03985_),
    .C(_03986_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08912_ (.I(_03855_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(\stack[10][7] ),
    .A2(_03976_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08914_ (.A1(_03887_),
    .A2(_03984_),
    .B1(_03969_),
    .B2(_03987_),
    .C(_03988_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08915_ (.I(_03669_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08916_ (.A1(_01605_),
    .A2(_03771_),
    .A3(_03821_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08917_ (.I(_03990_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08918_ (.A1(_03989_),
    .A2(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08919_ (.I(_03187_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08920_ (.I(_01690_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08921_ (.A1(_03827_),
    .A2(_03993_),
    .A3(_03994_),
    .A4(_03675_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08922_ (.I(_03678_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08923_ (.A1(_03996_),
    .A2(_03991_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08924_ (.A1(_03973_),
    .A2(_03995_),
    .A3(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08925_ (.I(_03998_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08926_ (.A1(\stack[13][0] ),
    .A2(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08927_ (.I(_03995_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08928_ (.A1(_03898_),
    .A2(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08929_ (.A1(_03890_),
    .A2(_03992_),
    .B(_04000_),
    .C(_04002_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08930_ (.I(_03992_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08931_ (.I(_01792_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08932_ (.A1(_04004_),
    .A2(_04001_),
    .B1(_03999_),
    .B2(\stack[13][1] ),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08933_ (.A1(_03952_),
    .A2(_04003_),
    .B(_04005_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08934_ (.I(_01824_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08935_ (.A1(_04006_),
    .A2(_04001_),
    .B1(_03999_),
    .B2(\stack[13][2] ),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08936_ (.A1(_03954_),
    .A2(_04003_),
    .B(_04007_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08937_ (.I(_01856_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08938_ (.I(_03998_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08939_ (.A1(_04008_),
    .A2(_04001_),
    .B1(_04009_),
    .B2(\stack[13][3] ),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08940_ (.A1(_03957_),
    .A2(_04003_),
    .B(_04010_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08941_ (.I(_01887_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08942_ (.A1(_04011_),
    .A2(_03995_),
    .B1(_04009_),
    .B2(\stack[13][4] ),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08943_ (.A1(_03959_),
    .A2(_04003_),
    .B(_04012_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_01922_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08945_ (.A1(_04013_),
    .A2(_03995_),
    .B1(_04009_),
    .B2(\stack[13][5] ),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08946_ (.A1(_03961_),
    .A2(_03992_),
    .B(_04014_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08947_ (.I(_03691_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08948_ (.A1(_03230_),
    .A2(_03848_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(_04015_),
    .A2(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08950_ (.A1(_03851_),
    .A2(_03997_),
    .B1(_04009_),
    .B2(\stack[13][6] ),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08951_ (.A1(_03846_),
    .A2(_04017_),
    .B(_04018_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08952_ (.I(_03853_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08953_ (.A1(\stack[13][7] ),
    .A2(_03999_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08954_ (.A1(_04019_),
    .A2(_04017_),
    .B1(_03992_),
    .B2(_03987_),
    .C(_04020_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08955_ (.A1(_01617_),
    .A2(_03201_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08956_ (.I(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08957_ (.I(_04022_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08958_ (.I(_01757_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08959_ (.I(_01684_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08960_ (.I(_01691_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08961_ (.A1(_03186_),
    .A2(_04025_),
    .A3(_04026_),
    .A4(_03234_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08962_ (.I(_04027_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08963_ (.A1(_03973_),
    .A2(_04027_),
    .A3(_04021_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08964_ (.I(_04029_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08965_ (.A1(_04024_),
    .A2(_04028_),
    .B1(_04030_),
    .B2(\stack[0][0] ),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08966_ (.A1(_03819_),
    .A2(_04023_),
    .B(_04031_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08967_ (.A1(_04004_),
    .A2(_04028_),
    .B1(_04030_),
    .B2(\stack[0][1] ),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03952_),
    .A2(_04023_),
    .B(_04032_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08969_ (.A1(_04006_),
    .A2(_04028_),
    .B1(_04030_),
    .B2(\stack[0][2] ),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08970_ (.A1(_03954_),
    .A2(_04023_),
    .B(_04033_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08971_ (.A1(_04008_),
    .A2(_04028_),
    .B1(_04030_),
    .B2(\stack[0][3] ),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08972_ (.A1(_03957_),
    .A2(_04023_),
    .B(_04034_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08973_ (.I(_04029_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08974_ (.A1(_04011_),
    .A2(_04027_),
    .B1(_04035_),
    .B2(\stack[0][4] ),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08975_ (.A1(_03959_),
    .A2(_04022_),
    .B(_04036_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08976_ (.A1(_04013_),
    .A2(_04027_),
    .B1(_04035_),
    .B2(\stack[0][5] ),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08977_ (.A1(_03961_),
    .A2(_04022_),
    .B(_04037_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08978_ (.I(_03731_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08979_ (.A1(_01932_),
    .A2(_03235_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08980_ (.I(_03237_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08981_ (.A1(_04040_),
    .A2(_04021_),
    .B1(_04035_),
    .B2(\stack[0][6] ),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_04038_),
    .A2(_04039_),
    .B(_04041_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08983_ (.A1(_03937_),
    .A2(_04021_),
    .B1(_04035_),
    .B2(\stack[0][7] ),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08984_ (.A1(_03936_),
    .A2(_04039_),
    .B(_04042_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08985_ (.A1(_03672_),
    .A2(_03993_),
    .A3(_03944_),
    .A4(_03675_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08986_ (.A1(_03679_),
    .A2(_03939_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08987_ (.A1(_03973_),
    .A2(_04043_),
    .A3(_04044_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08988_ (.I(_04045_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(\stack[25][0] ),
    .A2(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08990_ (.I(_04043_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08991_ (.A1(_03918_),
    .A2(_04048_),
    .B1(_04044_),
    .B2(_03866_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08992_ (.A1(_04047_),
    .A2(_04049_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08993_ (.I(_03868_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08994_ (.A1(_03669_),
    .A2(_03941_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08995_ (.I(_04051_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08996_ (.A1(_04004_),
    .A2(_04048_),
    .B1(_04046_),
    .B2(\stack[25][1] ),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08997_ (.A1(_04050_),
    .A2(_04052_),
    .B(_04053_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08998_ (.I(_03712_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08999_ (.A1(_04006_),
    .A2(_04048_),
    .B1(_04046_),
    .B2(\stack[25][2] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09000_ (.A1(_04054_),
    .A2(_04052_),
    .B(_04055_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09001_ (.I(_03716_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09002_ (.I(_04045_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09003_ (.A1(_04008_),
    .A2(_04048_),
    .B1(_04057_),
    .B2(\stack[25][3] ),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09004_ (.A1(_04056_),
    .A2(_04052_),
    .B(_04058_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09005_ (.I(_01860_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09006_ (.A1(_04011_),
    .A2(_04043_),
    .B1(_04057_),
    .B2(\stack[25][4] ),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09007_ (.A1(_04059_),
    .A2(_04052_),
    .B(_04060_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09008_ (.I(_01892_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09009_ (.A1(_04013_),
    .A2(_04043_),
    .B1(_04057_),
    .B2(\stack[25][5] ),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09010_ (.A1(_04061_),
    .A2(_04051_),
    .B(_04062_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(_04015_),
    .A2(_03964_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09012_ (.A1(_04040_),
    .A2(_04044_),
    .B1(_04057_),
    .B2(\stack[25][6] ),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09013_ (.A1(_04038_),
    .A2(_04063_),
    .B(_04064_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09014_ (.A1(\stack[25][7] ),
    .A2(_04046_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09015_ (.A1(_04019_),
    .A2(_04063_),
    .B1(_04051_),
    .B2(_03987_),
    .C(_04065_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09016_ (.I(_03889_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09017_ (.A1(_03989_),
    .A2(_03824_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09018_ (.I(_04067_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09019_ (.A1(_03827_),
    .A2(_03993_),
    .A3(_03944_),
    .A4(_03675_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09020_ (.I(_04069_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09021_ (.I(_03780_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09022_ (.A1(_03996_),
    .A2(_03822_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09023_ (.A1(_04071_),
    .A2(_04069_),
    .A3(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09024_ (.I(_04073_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09025_ (.A1(_04024_),
    .A2(_04070_),
    .B1(_04074_),
    .B2(\stack[9][0] ),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_04066_),
    .A2(_04068_),
    .B(_04075_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09027_ (.A1(_04004_),
    .A2(_04070_),
    .B1(_04074_),
    .B2(\stack[9][1] ),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09028_ (.A1(_04050_),
    .A2(_04068_),
    .B(_04076_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09029_ (.A1(_04006_),
    .A2(_04070_),
    .B1(_04074_),
    .B2(\stack[9][2] ),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09030_ (.A1(_04054_),
    .A2(_04068_),
    .B(_04077_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09031_ (.I(_04073_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09032_ (.A1(_04008_),
    .A2(_04070_),
    .B1(_04078_),
    .B2(\stack[9][3] ),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09033_ (.A1(_04056_),
    .A2(_04068_),
    .B(_04079_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09034_ (.A1(_04011_),
    .A2(_04069_),
    .B1(_04078_),
    .B2(\stack[9][4] ),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09035_ (.A1(_04059_),
    .A2(_04067_),
    .B(_04080_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09036_ (.A1(_04013_),
    .A2(_04069_),
    .B1(_04078_),
    .B2(\stack[9][5] ),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09037_ (.A1(_04061_),
    .A2(_04067_),
    .B(_04081_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(_04015_),
    .A2(_03849_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09039_ (.A1(_04040_),
    .A2(_04072_),
    .B1(_04078_),
    .B2(\stack[9][6] ),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_04038_),
    .A2(_04082_),
    .B(_04083_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09041_ (.A1(\stack[9][7] ),
    .A2(_04074_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09042_ (.A1(_04019_),
    .A2(_04082_),
    .B1(_04067_),
    .B2(_03987_),
    .C(_04084_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09043_ (.A1(_03636_),
    .A2(_01685_),
    .A3(_01930_),
    .A4(_03663_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09044_ (.A1(_03629_),
    .A2(_03770_),
    .A3(_01616_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09045_ (.I(_04086_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_03743_),
    .A2(_04087_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09047_ (.A1(_03740_),
    .A2(_04085_),
    .A3(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09048_ (.I(_04089_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09049_ (.A1(\stack[23][0] ),
    .A2(_04090_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09050_ (.I(_04085_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09051_ (.I(_04088_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09052_ (.A1(_03918_),
    .A2(_04092_),
    .B1(_04093_),
    .B2(_03866_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_04091_),
    .A2(_04094_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09054_ (.A1(_03870_),
    .A2(_04087_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09055_ (.I(_04089_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(\stack[23][1] ),
    .A2(_04096_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(_03752_),
    .A2(_04092_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09058_ (.A1(_03869_),
    .A2(_04095_),
    .B(_04097_),
    .C(_04098_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09059_ (.A1(\stack[23][2] ),
    .A2(_04090_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09060_ (.I(_00919_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09061_ (.A1(_03755_),
    .A2(_04092_),
    .B1(_04093_),
    .B2(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09062_ (.A1(_04099_),
    .A2(_04101_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(\stack[23][3] ),
    .A2(_04090_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09064_ (.I(_00983_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09065_ (.A1(_03758_),
    .A2(_04085_),
    .B1(_04093_),
    .B2(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(_04102_),
    .A2(_04104_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(\stack[23][4] ),
    .A2(_04096_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(_03762_),
    .A2(_04092_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09069_ (.A1(_03879_),
    .A2(_04095_),
    .B(_04105_),
    .C(_04106_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09070_ (.A1(_03228_),
    .A2(_04085_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(\stack[23][5] ),
    .A2(_04090_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09072_ (.A1(_03882_),
    .A2(_04095_),
    .B(_04107_),
    .C(_04108_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09073_ (.A1(_03230_),
    .A2(_03661_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_03663_),
    .A2(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09075_ (.A1(_04040_),
    .A2(_04093_),
    .B1(_04096_),
    .B2(\stack[23][6] ),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09076_ (.A1(_04038_),
    .A2(_04110_),
    .B(_04111_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09077_ (.I(_03855_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(\stack[23][7] ),
    .A2(_04096_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09079_ (.A1(_04019_),
    .A2(_04110_),
    .B1(_04095_),
    .B2(_04112_),
    .C(_04113_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09080_ (.A1(_03820_),
    .A2(_03941_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09081_ (.I(_04114_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09082_ (.A1(_03672_),
    .A2(_03993_),
    .A3(_01929_),
    .A4(_03192_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09083_ (.I(_04116_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09084_ (.A1(_03820_),
    .A2(_03940_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09085_ (.A1(_04071_),
    .A2(_04116_),
    .A3(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09086_ (.I(_04119_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09087_ (.A1(_04024_),
    .A2(_04117_),
    .B1(_04120_),
    .B2(\stack[24][0] ),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09088_ (.A1(_04066_),
    .A2(_04115_),
    .B(_04121_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09089_ (.I(_01792_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09090_ (.A1(_04122_),
    .A2(_04117_),
    .B1(_04120_),
    .B2(\stack[24][1] ),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09091_ (.A1(_04050_),
    .A2(_04115_),
    .B(_04123_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09092_ (.I(_01824_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09093_ (.A1(_04124_),
    .A2(_04117_),
    .B1(_04120_),
    .B2(\stack[24][2] ),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_04054_),
    .A2(_04115_),
    .B(_04125_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09095_ (.I(_01856_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09096_ (.I(_04119_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09097_ (.A1(_04126_),
    .A2(_04117_),
    .B1(_04127_),
    .B2(\stack[24][3] ),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09098_ (.A1(_04056_),
    .A2(_04115_),
    .B(_04128_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09099_ (.I(_01887_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09100_ (.A1(_04129_),
    .A2(_04116_),
    .B1(_04127_),
    .B2(\stack[24][4] ),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09101_ (.A1(_04059_),
    .A2(_04114_),
    .B(_04130_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09102_ (.I(_01922_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09103_ (.A1(_04131_),
    .A2(_04116_),
    .B1(_04127_),
    .B2(\stack[24][5] ),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09104_ (.A1(_04061_),
    .A2(_04114_),
    .B(_04132_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09105_ (.I(_03731_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(_03847_),
    .A2(_03964_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09107_ (.I(_01124_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09108_ (.A1(_04135_),
    .A2(_04118_),
    .B1(_04127_),
    .B2(\stack[24][6] ),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09109_ (.A1(_04133_),
    .A2(_04134_),
    .B(_04136_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09110_ (.I(_03853_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(\stack[24][7] ),
    .A2(_04120_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09112_ (.A1(_04137_),
    .A2(_04134_),
    .B1(_04114_),
    .B2(_04112_),
    .C(_04138_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09113_ (.A1(net42),
    .A2(net67),
    .A3(_01626_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09114_ (.I(_04139_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09115_ (.I(_04140_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09116_ (.A1(_03282_),
    .A2(_04141_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09117_ (.A1(_01638_),
    .A2(_03643_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09118_ (.I(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09119_ (.I(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09120_ (.I(_03635_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09121_ (.A1(_04145_),
    .A2(_04025_),
    .A3(_04026_),
    .A4(_01712_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09122_ (.I(_04146_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09123_ (.A1(_04071_),
    .A2(_04146_),
    .A3(_04142_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09124_ (.I(_04148_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09125_ (.A1(_04024_),
    .A2(_04147_),
    .B1(_04149_),
    .B2(\stack[18][0] ),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_04066_),
    .A2(_04144_),
    .B(_04150_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09127_ (.A1(_04122_),
    .A2(_04147_),
    .B1(_04149_),
    .B2(\stack[18][1] ),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09128_ (.A1(_04050_),
    .A2(_04144_),
    .B(_04151_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09129_ (.A1(_04124_),
    .A2(_04147_),
    .B1(_04149_),
    .B2(\stack[18][2] ),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09130_ (.A1(_04054_),
    .A2(_04144_),
    .B(_04152_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09131_ (.I(_04148_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09132_ (.A1(_04126_),
    .A2(_04147_),
    .B1(_04153_),
    .B2(\stack[18][3] ),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09133_ (.A1(_04056_),
    .A2(_04144_),
    .B(_04154_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09134_ (.A1(_04129_),
    .A2(_04146_),
    .B1(_04153_),
    .B2(\stack[18][4] ),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09135_ (.A1(_04059_),
    .A2(_04143_),
    .B(_04155_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09136_ (.A1(_04131_),
    .A2(_04146_),
    .B1(_04153_),
    .B2(\stack[18][5] ),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09137_ (.A1(_04061_),
    .A2(_04143_),
    .B(_04156_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(_03909_),
    .A2(_03662_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09139_ (.A1(\stack[18][6] ),
    .A2(_04149_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09140_ (.A1(_03238_),
    .A2(_04142_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09141_ (.A1(_03963_),
    .A2(_04157_),
    .B(_04158_),
    .C(_04159_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09142_ (.A1(_03937_),
    .A2(_04142_),
    .B1(_04153_),
    .B2(\stack[18][7] ),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09143_ (.A1(_03936_),
    .A2(_04157_),
    .B(_04160_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09144_ (.A1(_03186_),
    .A2(_04025_),
    .A3(_04026_),
    .A4(_03691_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09145_ (.A1(_01617_),
    .A2(_03679_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09146_ (.A1(_04071_),
    .A2(_04161_),
    .A3(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09147_ (.I(_04163_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(\stack[1][0] ),
    .A2(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09149_ (.I(_04161_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09150_ (.I(_00842_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09151_ (.A1(_03918_),
    .A2(_04166_),
    .B1(_04162_),
    .B2(_04167_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09152_ (.A1(_04165_),
    .A2(_04168_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09153_ (.I(_03868_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09154_ (.A1(_01618_),
    .A2(_03989_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09155_ (.I(_04170_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09156_ (.A1(_04122_),
    .A2(_04166_),
    .B1(_04164_),
    .B2(\stack[1][1] ),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09157_ (.A1(_04169_),
    .A2(_04171_),
    .B(_04172_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09158_ (.I(_03712_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09159_ (.A1(_04124_),
    .A2(_04166_),
    .B1(_04164_),
    .B2(\stack[1][2] ),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_04173_),
    .A2(_04171_),
    .B(_04174_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09161_ (.I(_03716_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09162_ (.A1(_04126_),
    .A2(_04166_),
    .B1(_04164_),
    .B2(\stack[1][3] ),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09163_ (.A1(_04175_),
    .A2(_04171_),
    .B(_04176_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09164_ (.I(_03721_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09165_ (.I(_04163_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09166_ (.A1(_04129_),
    .A2(_04161_),
    .B1(_04178_),
    .B2(\stack[1][4] ),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09167_ (.A1(_04177_),
    .A2(_04171_),
    .B(_04179_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09168_ (.I(_03728_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09169_ (.A1(_04131_),
    .A2(_04161_),
    .B1(_04178_),
    .B2(\stack[1][5] ),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09170_ (.A1(_04180_),
    .A2(_04170_),
    .B(_04181_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(_01932_),
    .A2(_03692_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09172_ (.A1(_04135_),
    .A2(_04162_),
    .B1(_04178_),
    .B2(\stack[1][6] ),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09173_ (.A1(_04133_),
    .A2(_04182_),
    .B(_04183_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09174_ (.A1(_03937_),
    .A2(_04162_),
    .B1(_04178_),
    .B2(\stack[1][7] ),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09175_ (.A1(_03936_),
    .A2(_04182_),
    .B(_04184_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09176_ (.I(_03780_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09177_ (.A1(_04145_),
    .A2(_04025_),
    .A3(_03777_),
    .A4(_03233_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09178_ (.A1(_03202_),
    .A2(_04086_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09179_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09180_ (.I(_04188_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09181_ (.A1(\stack[20][0] ),
    .A2(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09182_ (.I(_03207_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09183_ (.I(_04186_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09184_ (.I(_04187_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09185_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_04193_),
    .B2(_04167_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_04190_),
    .A2(_04194_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09187_ (.I(_04193_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09188_ (.I(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09189_ (.A1(_04122_),
    .A2(_04192_),
    .B1(_04189_),
    .B2(\stack[20][1] ),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09190_ (.A1(_04169_),
    .A2(_04196_),
    .B(_04197_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09191_ (.A1(_04124_),
    .A2(_04192_),
    .B1(_04189_),
    .B2(\stack[20][2] ),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09192_ (.A1(_04173_),
    .A2(_04196_),
    .B(_04198_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09193_ (.A1(_04126_),
    .A2(_04192_),
    .B1(_04189_),
    .B2(\stack[20][3] ),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_04175_),
    .A2(_04196_),
    .B(_04199_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09195_ (.I(_04188_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09196_ (.A1(_04129_),
    .A2(_04186_),
    .B1(_04200_),
    .B2(\stack[20][4] ),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09197_ (.A1(_04177_),
    .A2(_04196_),
    .B(_04201_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09198_ (.A1(_04131_),
    .A2(_04186_),
    .B1(_04200_),
    .B2(\stack[20][5] ),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09199_ (.A1(_04180_),
    .A2(_04195_),
    .B(_04202_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_03235_),
    .A2(_04109_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09201_ (.A1(_04135_),
    .A2(_04193_),
    .B1(_04200_),
    .B2(\stack[20][6] ),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09202_ (.A1(_04133_),
    .A2(_04203_),
    .B(_04204_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09203_ (.I(_01990_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09204_ (.I(_01170_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09205_ (.A1(_04206_),
    .A2(_04193_),
    .B1(_04200_),
    .B2(\stack[20][7] ),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09206_ (.A1(_04205_),
    .A2(_04203_),
    .B(_04207_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09207_ (.A1(_03989_),
    .A2(_04087_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09208_ (.I(_03187_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09209_ (.A1(_04145_),
    .A2(_04209_),
    .A3(_03777_),
    .A4(_03690_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09210_ (.A1(_03996_),
    .A2(_04087_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09211_ (.A1(_04185_),
    .A2(_04210_),
    .A3(_04211_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09212_ (.I(_04212_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09213_ (.A1(\stack[21][0] ),
    .A2(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09214_ (.I(_04210_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_03898_),
    .A2(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09216_ (.A1(_01182_),
    .A2(_04208_),
    .B(_04214_),
    .C(_04216_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09217_ (.I(_04208_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09218_ (.I(_01792_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09219_ (.A1(_04218_),
    .A2(_04215_),
    .B1(_04213_),
    .B2(\stack[21][1] ),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09220_ (.A1(_04169_),
    .A2(_04217_),
    .B(_04219_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09221_ (.I(_01824_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09222_ (.A1(_04220_),
    .A2(_04215_),
    .B1(_04213_),
    .B2(\stack[21][2] ),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09223_ (.A1(_04173_),
    .A2(_04217_),
    .B(_04221_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09224_ (.I(_01856_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09225_ (.I(_04212_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09226_ (.A1(_04222_),
    .A2(_04215_),
    .B1(_04223_),
    .B2(\stack[21][3] ),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09227_ (.A1(_04175_),
    .A2(_04217_),
    .B(_04224_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09228_ (.I(_01887_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09229_ (.A1(_04225_),
    .A2(_04210_),
    .B1(_04223_),
    .B2(\stack[21][4] ),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_04177_),
    .A2(_04217_),
    .B(_04226_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09231_ (.I(_01922_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09232_ (.A1(_04227_),
    .A2(_04210_),
    .B1(_04223_),
    .B2(\stack[21][5] ),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09233_ (.A1(_04180_),
    .A2(_04208_),
    .B(_04228_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_04015_),
    .A2(_04109_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09235_ (.A1(_04135_),
    .A2(_04211_),
    .B1(_04223_),
    .B2(\stack[21][6] ),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09236_ (.A1(_04133_),
    .A2(_04229_),
    .B(_04230_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(\stack[21][7] ),
    .A2(_04213_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09238_ (.A1(_04137_),
    .A2(_04229_),
    .B1(_04208_),
    .B2(_04112_),
    .C(_04231_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09239_ (.A1(_01715_),
    .A2(_04086_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09240_ (.I(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09241_ (.I(_04233_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09242_ (.A1(_04145_),
    .A2(_04209_),
    .A3(_03828_),
    .A4(_01712_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09243_ (.I(_04235_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09244_ (.A1(_04185_),
    .A2(_04235_),
    .A3(_04232_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09245_ (.I(_04237_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09246_ (.A1(_01758_),
    .A2(_04236_),
    .B1(_04238_),
    .B2(\stack[22][0] ),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09247_ (.A1(_04066_),
    .A2(_04234_),
    .B(_04239_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09248_ (.A1(_04218_),
    .A2(_04236_),
    .B1(_04238_),
    .B2(\stack[22][1] ),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09249_ (.A1(_04169_),
    .A2(_04234_),
    .B(_04240_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09250_ (.A1(_04220_),
    .A2(_04236_),
    .B1(_04238_),
    .B2(\stack[22][2] ),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09251_ (.A1(_04173_),
    .A2(_04234_),
    .B(_04241_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09252_ (.I(_04237_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09253_ (.A1(_04222_),
    .A2(_04236_),
    .B1(_04242_),
    .B2(\stack[22][3] ),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09254_ (.A1(_04175_),
    .A2(_04234_),
    .B(_04243_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09255_ (.A1(_04225_),
    .A2(_04235_),
    .B1(_04242_),
    .B2(\stack[22][4] ),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09256_ (.A1(_04177_),
    .A2(_04233_),
    .B(_04244_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09257_ (.A1(_04227_),
    .A2(_04235_),
    .B1(_04242_),
    .B2(\stack[22][5] ),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09258_ (.A1(_04180_),
    .A2(_04233_),
    .B(_04245_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09259_ (.A1(_03909_),
    .A2(_04109_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(\stack[22][6] ),
    .A2(_04238_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09261_ (.A1(_03908_),
    .A2(_04246_),
    .B1(_04233_),
    .B2(_03733_),
    .C(_04247_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09262_ (.A1(_04206_),
    .A2(_04232_),
    .B1(_04242_),
    .B2(\stack[22][7] ),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09263_ (.A1(_04205_),
    .A2(_04246_),
    .B(_04248_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09264_ (.I(net143),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09265_ (.I(_04249_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09266_ (.I(net256),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09267_ (.I(net141),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09268_ (.A1(net77),
    .A2(net193),
    .B(\mem.dff_data_ready ),
    .C(\mem.io_data_ready ),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09269_ (.A1(_01171_),
    .A2(_04253_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09270_ (.A1(_04250_),
    .A2(_04251_),
    .A3(_04252_),
    .A4(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09271_ (.I(_04252_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09272_ (.A1(net256),
    .A2(_04256_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(_04249_),
    .A2(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09274_ (.A1(_03620_),
    .A2(_04258_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09275_ (.A1(_01662_),
    .A2(_01663_),
    .A3(_01664_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09276_ (.I(_04260_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09277_ (.A1(_01661_),
    .A2(_04259_),
    .A3(_04261_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09278_ (.A1(_03621_),
    .A2(_04255_),
    .B(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09279_ (.I(_04263_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09280_ (.I(_04264_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09281_ (.I(_03622_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09282_ (.I(_03241_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09283_ (.I(_01172_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09284_ (.A1(net78),
    .A2(_02289_),
    .B1(_00760_),
    .B2(net94),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09285_ (.I(\mem.sram_enable ),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09286_ (.A1(net85),
    .A2(_00761_),
    .B1(_00762_),
    .B2(net108),
    .C(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09287_ (.A1(_04269_),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09288_ (.A1(_04268_),
    .A2(\mem.dff_data_out[0] ),
    .B(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09289_ (.I(_03241_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09290_ (.A1(\mem.io_data_out[0] ),
    .A2(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09291_ (.A1(_04267_),
    .A2(_04273_),
    .B(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09292_ (.A1(_03622_),
    .A2(_01727_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09293_ (.A1(_04266_),
    .A2(_04276_),
    .B(_04277_),
    .C(_04264_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09294_ (.A1(_01212_),
    .A2(_04265_),
    .B(_04278_),
    .C(_03627_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09295_ (.A1(net95),
    .A2(net230),
    .B1(net229),
    .B2(net86),
    .C1(net228),
    .C2(net109),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_03099_),
    .A2(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09297_ (.I(_04270_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09298_ (.A1(net89),
    .A2(_03099_),
    .B(_04280_),
    .C(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09299_ (.I(_04268_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09300_ (.A1(_04283_),
    .A2(\mem.dff_data_out[1] ),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09301_ (.A1(_04282_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09302_ (.I0(\mem.io_data_out[1] ),
    .I1(_04285_),
    .S(_03242_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09303_ (.A1(_04266_),
    .A2(_04286_),
    .B(_04263_),
    .C(_03624_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09304_ (.I(_02003_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09305_ (.I(_04288_),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09306_ (.A1(_01196_),
    .A2(_04265_),
    .B(_04287_),
    .C(_04289_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09307_ (.A1(net100),
    .A2(_02289_),
    .B1(_00760_),
    .B2(net96),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09308_ (.I(_00761_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09309_ (.I(_00762_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09310_ (.A1(net87),
    .A2(_04291_),
    .B1(_04292_),
    .B2(net79),
    .C(_04270_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09311_ (.A1(_04290_),
    .A2(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09312_ (.A1(_04268_),
    .A2(\mem.dff_data_out[2] ),
    .B(_04294_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09313_ (.A1(\mem.io_data_out[2] ),
    .A2(_04274_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09314_ (.A1(_04267_),
    .A2(_04295_),
    .B(_04296_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09315_ (.I(_03621_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09316_ (.I(_01800_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09317_ (.A1(_04298_),
    .A2(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09318_ (.I(_04263_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09319_ (.A1(_04266_),
    .A2(_04297_),
    .B(_04300_),
    .C(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09320_ (.A1(_01207_),
    .A2(_04265_),
    .B(_04302_),
    .C(_04289_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09321_ (.I(_03622_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09322_ (.I(_00758_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09323_ (.A1(net103),
    .A2(_04304_),
    .B1(_02134_),
    .B2(net97),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09324_ (.I(_04270_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09325_ (.A1(net88),
    .A2(_04291_),
    .B1(_04292_),
    .B2(net80),
    .C(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09326_ (.A1(_04305_),
    .A2(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09327_ (.A1(_04268_),
    .A2(\mem.dff_data_out[3] ),
    .B(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09328_ (.A1(\mem.io_data_out[3] ),
    .A2(_04274_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09329_ (.A1(_04267_),
    .A2(_04309_),
    .B(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09330_ (.I(_01833_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09331_ (.A1(_04298_),
    .A2(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09332_ (.A1(_04303_),
    .A2(_04311_),
    .B(_04313_),
    .C(_04301_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09333_ (.A1(_01227_),
    .A2(_04265_),
    .B(_04314_),
    .C(_04289_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09334_ (.I(_04264_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09335_ (.A1(net104),
    .A2(_04304_),
    .B1(_02618_),
    .B2(net98),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09336_ (.A1(net90),
    .A2(_03042_),
    .B1(_03014_),
    .B2(net81),
    .C(_04306_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09337_ (.A1(_04316_),
    .A2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09338_ (.A1(_04283_),
    .A2(\mem.dff_data_out[4] ),
    .B(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09339_ (.I(_03241_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09340_ (.A1(\mem.io_data_out[4] ),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09341_ (.A1(_03242_),
    .A2(_04319_),
    .B(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09342_ (.I(_03620_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09343_ (.I(_04323_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09344_ (.I(_01864_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09345_ (.A1(_04324_),
    .A2(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09346_ (.A1(_04303_),
    .A2(_04322_),
    .B(_04326_),
    .C(_04301_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09347_ (.A1(_01186_),
    .A2(_04315_),
    .B(_04327_),
    .C(_04289_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09348_ (.A1(net105),
    .A2(_04304_),
    .B1(_02134_),
    .B2(net99),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09349_ (.A1(net91),
    .A2(_04291_),
    .B1(_04292_),
    .B2(net82),
    .C(_04306_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09350_ (.A1(_04328_),
    .A2(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09351_ (.A1(_04283_),
    .A2(\mem.dff_data_out[5] ),
    .B(_04330_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09352_ (.A1(\mem.io_data_out[5] ),
    .A2(_04320_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09353_ (.A1(_04320_),
    .A2(_04331_),
    .B(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09354_ (.A1(_04298_),
    .A2(_01896_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09355_ (.A1(_04303_),
    .A2(_04333_),
    .B(_04334_),
    .C(_04301_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09356_ (.I(_02003_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09357_ (.I(_04336_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09358_ (.A1(_01214_),
    .A2(_04315_),
    .B(_04335_),
    .C(_04337_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09359_ (.A1(_01723_),
    .A2(_01628_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09360_ (.I(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09361_ (.A1(net106),
    .A2(_04304_),
    .B1(_02134_),
    .B2(net101),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09362_ (.A1(net92),
    .A2(_04291_),
    .B1(_04292_),
    .B2(net83),
    .C(_04306_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09363_ (.A1(_01172_),
    .A2(\mem.dff_data_out[6] ),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09364_ (.A1(_04340_),
    .A2(_04341_),
    .B(_04342_),
    .C(_04274_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09365_ (.A1(\mem.io_data_out[6] ),
    .A2(_04267_),
    .B(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09366_ (.A1(_04339_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09367_ (.A1(_04324_),
    .A2(_01960_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09368_ (.A1(_04264_),
    .A2(_04345_),
    .A3(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09369_ (.A1(_01218_),
    .A2(_04315_),
    .B(_04347_),
    .C(_04337_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09370_ (.A1(net107),
    .A2(_03099_),
    .B1(_02618_),
    .B2(net102),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09371_ (.A1(net93),
    .A2(_03042_),
    .B1(_03014_),
    .B2(net84),
    .C(_04281_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09372_ (.A1(_04348_),
    .A2(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09373_ (.A1(_04283_),
    .A2(\mem.dff_data_out[7] ),
    .B(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09374_ (.A1(\mem.io_data_out[7] ),
    .A2(_04320_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09375_ (.A1(_03242_),
    .A2(_04351_),
    .B(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09376_ (.I(_01765_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09377_ (.A1(_04354_),
    .A2(_01986_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09378_ (.A1(_04354_),
    .A2(net64),
    .B(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09379_ (.A1(_04298_),
    .A2(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09380_ (.A1(_04303_),
    .A2(_04353_),
    .B(_04357_),
    .C(_04263_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09381_ (.A1(_01222_),
    .A2(_04315_),
    .B(_04358_),
    .C(_04337_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09382_ (.I(net128),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09383_ (.A1(_01630_),
    .A2(_03616_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09384_ (.A1(_01659_),
    .A2(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09385_ (.I(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09386_ (.A1(_04261_),
    .A2(_04362_),
    .B(_03625_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09387_ (.I(_04363_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09388_ (.I(_04364_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09389_ (.A1(_04277_),
    .A2(_04364_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09390_ (.A1(_01198_),
    .A2(_01200_),
    .A3(_01202_),
    .B(_01575_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09391_ (.I(_04367_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09392_ (.I(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09393_ (.A1(\exec.out_of_order_exec ),
    .A2(_04359_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09394_ (.I(_04367_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09395_ (.A1(_03889_),
    .A2(_04371_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09396_ (.A1(_04369_),
    .A2(_04370_),
    .B(_04372_),
    .C(_04266_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09397_ (.I(_01644_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09398_ (.I(_04374_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09399_ (.A1(_04359_),
    .A2(_04365_),
    .B1(_04366_),
    .B2(_04373_),
    .C(_04375_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09400_ (.I(net139),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09401_ (.I(_04376_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09402_ (.A1(\exec.out_of_order_exec ),
    .A2(_04359_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09403_ (.A1(_04376_),
    .A2(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09404_ (.I(_04367_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09405_ (.A1(_01762_),
    .A2(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09406_ (.I(_04323_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09407_ (.A1(_04369_),
    .A2(_04379_),
    .B(_04381_),
    .C(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09408_ (.I(_04364_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09409_ (.A1(_03624_),
    .A2(_04384_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09410_ (.A1(_04377_),
    .A2(_04365_),
    .B1(_04383_),
    .B2(_04385_),
    .C(_04375_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09411_ (.I(net257),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09412_ (.I(_04338_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09413_ (.I(_04387_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09414_ (.A1(net257),
    .A2(net139),
    .A3(_04378_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(net139),
    .A2(_04378_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09416_ (.A1(_04386_),
    .A2(_04390_),
    .B(_04367_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09417_ (.A1(_00919_),
    .A2(_04368_),
    .B1(_04389_),
    .B2(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09418_ (.A1(_04388_),
    .A2(_04392_),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09419_ (.A1(_04300_),
    .A2(_04384_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09420_ (.A1(_04386_),
    .A2(_04365_),
    .B1(_04393_),
    .B2(_04394_),
    .C(_04375_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09421_ (.I(net153),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09422_ (.A1(_04395_),
    .A2(_04389_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(_01827_),
    .A2(_04380_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09424_ (.A1(_04369_),
    .A2(_04396_),
    .B(_04397_),
    .C(_04382_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09425_ (.I(_04363_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09426_ (.A1(_04313_),
    .A2(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09427_ (.I(_04374_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09428_ (.A1(_04395_),
    .A2(_04365_),
    .B1(_04398_),
    .B2(_04400_),
    .C(_04401_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09429_ (.I(_03621_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09430_ (.I(_04402_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09431_ (.A1(_04395_),
    .A2(_04389_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09432_ (.A1(net154),
    .A2(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09433_ (.I(net154),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09434_ (.A1(_04406_),
    .A2(_04404_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(_01027_),
    .A2(_04368_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09436_ (.A1(_04371_),
    .A2(_04405_),
    .A3(_04407_),
    .B(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09437_ (.A1(_04403_),
    .A2(_04409_),
    .B(_04399_),
    .C(_04326_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09438_ (.I(_04260_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09439_ (.I(_01624_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09440_ (.I(_04412_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(_04413_),
    .A2(_04323_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09442_ (.A1(_04411_),
    .A2(_04361_),
    .B(_04414_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09443_ (.A1(_04406_),
    .A2(_04415_),
    .B(_02000_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09444_ (.A1(_04410_),
    .A2(_04416_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09445_ (.I(net155),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09446_ (.I(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09447_ (.A1(_04417_),
    .A2(_04405_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(_01891_),
    .A2(_04380_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09449_ (.A1(_04369_),
    .A2(_04419_),
    .B(_04420_),
    .C(_04382_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09450_ (.A1(_04334_),
    .A2(_04399_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09451_ (.A1(_04418_),
    .A2(_04384_),
    .B1(_04421_),
    .B2(_04422_),
    .C(_04401_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09452_ (.I(net156),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(net155),
    .A2(_04405_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09454_ (.A1(_04423_),
    .A2(_04424_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(_01124_),
    .A2(_04368_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_04371_),
    .A2(_04425_),
    .B(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09457_ (.A1(_04403_),
    .A2(_04427_),
    .B(_04364_),
    .C(_04346_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09458_ (.I(_02009_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09459_ (.A1(_04423_),
    .A2(_04415_),
    .B(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09460_ (.A1(_04428_),
    .A2(_04430_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09461_ (.I(net157),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09462_ (.A1(net156),
    .A2(net155),
    .A3(_04405_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09463_ (.A1(_04431_),
    .A2(_04432_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09464_ (.A1(_03737_),
    .A2(_04380_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09465_ (.A1(_04371_),
    .A2(_04433_),
    .B(_04434_),
    .C(_04324_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09466_ (.A1(_04357_),
    .A2(_04399_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09467_ (.A1(_04431_),
    .A2(_04384_),
    .B1(_04435_),
    .B2(_04436_),
    .C(_04401_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09468_ (.A1(_01696_),
    .A2(_04411_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09469_ (.A1(_04338_),
    .A2(_01668_),
    .B1(_04360_),
    .B2(_04437_),
    .C(_03625_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09470_ (.I(_04438_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09471_ (.I(_04387_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09472_ (.I(_01667_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09473_ (.I(_01667_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09474_ (.A1(_01724_),
    .A2(net43),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09475_ (.A1(_01767_),
    .A2(_01725_),
    .B(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09476_ (.A1(_04442_),
    .A2(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09477_ (.A1(_01700_),
    .A2(_04441_),
    .B(_04445_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09478_ (.A1(_04440_),
    .A2(_04446_),
    .B(_04439_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_04403_),
    .A2(_03199_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09480_ (.A1(_01131_),
    .A2(_04439_),
    .B1(_04447_),
    .B2(_04448_),
    .C(_04401_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09481_ (.I(_04439_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09482_ (.A1(_01697_),
    .A2(_04261_),
    .B(_01668_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09483_ (.A1(_04402_),
    .A2(_04450_),
    .B(_04414_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_04442_),
    .A2(_01769_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09485_ (.A1(_01064_),
    .A2(_04441_),
    .B(_04452_),
    .C(_04339_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09486_ (.A1(_04440_),
    .A2(_03628_),
    .B(_04451_),
    .C(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_02000_),
    .A2(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09488_ (.A1(_01130_),
    .A2(_04449_),
    .B(_04455_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09489_ (.A1(_01667_),
    .A2(_04299_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09490_ (.A1(_04442_),
    .A2(_01595_),
    .B(_04456_),
    .C(_04387_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(_04388_),
    .A2(_01598_),
    .B(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09492_ (.A1(_04439_),
    .A2(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09493_ (.A1(_01286_),
    .A2(_04449_),
    .B(_04459_),
    .C(_04337_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09494_ (.A1(_04442_),
    .A2(_04312_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09495_ (.A1(_04441_),
    .A2(_01613_),
    .B(_04460_),
    .C(_04339_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09496_ (.A1(_04440_),
    .A2(_01615_),
    .B(_04451_),
    .C(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09497_ (.A1(_02000_),
    .A2(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09498_ (.A1(_00805_),
    .A2(_04449_),
    .B(_04463_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09499_ (.A1(_01661_),
    .A2(_01694_),
    .A3(_01257_),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09500_ (.A1(_04441_),
    .A2(_04325_),
    .B(_04464_),
    .C(_04402_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09501_ (.A1(_04382_),
    .A2(_01588_),
    .B(_04438_),
    .C(_04465_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09502_ (.I(_04336_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09503_ (.A1(_00850_),
    .A2(_04449_),
    .B(_04466_),
    .C(_04467_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09504_ (.I(_03281_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09505_ (.A1(_04468_),
    .A2(_03570_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09506_ (.A1(_01661_),
    .A2(_04259_),
    .A3(_04261_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09507_ (.A1(_03616_),
    .A2(_04444_),
    .A3(_04259_),
    .A4(_04437_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(\exec.out_of_order_exec ),
    .A2(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09509_ (.I(_02004_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09510_ (.A1(_04469_),
    .A2(_04471_),
    .B(_04472_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09511_ (.A1(_03616_),
    .A2(_04437_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09512_ (.A1(_04323_),
    .A2(_04473_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09513_ (.I(_04474_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09514_ (.A1(_04281_),
    .A2(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09515_ (.A1(_04299_),
    .A2(_04475_),
    .B(_04476_),
    .C(_04467_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09516_ (.A1(_04249_),
    .A2(_04251_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09517_ (.A1(_04249_),
    .A2(_01623_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09518_ (.A1(_04252_),
    .A2(_04478_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09519_ (.I(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09520_ (.A1(_04477_),
    .A2(_04480_),
    .B(_04402_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09521_ (.A1(_01171_),
    .A2(_04479_),
    .B(_04481_),
    .C(_04253_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09522_ (.A1(_01171_),
    .A2(_04481_),
    .B(_04482_),
    .C(_04467_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09523_ (.I(\cycles_per_ms[23] ),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09524_ (.I(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09525_ (.I(\delay_cycles[18] ),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09526_ (.I(\delay_cycles[15] ),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09527_ (.I(\delay_cycles[14] ),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09528_ (.I(\delay_cycles[13] ),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09529_ (.A1(\delay_cycles[3] ),
    .A2(\delay_cycles[2] ),
    .A3(\delay_cycles[1] ),
    .A4(\delay_cycles[0] ),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09530_ (.A1(\delay_cycles[6] ),
    .A2(\delay_cycles[5] ),
    .A3(\delay_cycles[4] ),
    .A4(_04489_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09531_ (.A1(\delay_cycles[9] ),
    .A2(\delay_cycles[8] ),
    .A3(\delay_cycles[7] ),
    .A4(_04490_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09532_ (.A1(\delay_cycles[12] ),
    .A2(\delay_cycles[11] ),
    .A3(\delay_cycles[10] ),
    .A4(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09533_ (.A1(_04486_),
    .A2(_04487_),
    .A3(_04488_),
    .A4(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09534_ (.A1(\delay_cycles[17] ),
    .A2(\delay_cycles[16] ),
    .A3(_04493_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09535_ (.I(_04494_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09536_ (.A1(\delay_cycles[19] ),
    .A2(_04485_),
    .A3(_04495_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09537_ (.A1(\delay_cycles[21] ),
    .A2(\delay_cycles[20] ),
    .A3(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09538_ (.A1(\delay_cycles[22] ),
    .A2(_04497_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09539_ (.A1(\delay_cycles[23] ),
    .A2(_04498_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09540_ (.I(\cycles_per_ms[22] ),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09541_ (.A1(\delay_cycles[22] ),
    .A2(_04497_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09542_ (.A1(\delay_cycles[20] ),
    .A2(_04496_),
    .B(\delay_cycles[21] ),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09543_ (.A1(_04497_),
    .A2(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09544_ (.I(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09545_ (.I(\cycles_per_ms[21] ),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09546_ (.A1(_04500_),
    .A2(_04501_),
    .B1(_04504_),
    .B2(_04505_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09547_ (.I(\cycles_per_ms[18] ),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09548_ (.A1(_04485_),
    .A2(_04495_),
    .Z(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09549_ (.I(\delay_cycles[16] ),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09550_ (.A1(\delay_cycles[18] ),
    .A2(\delay_cycles[17] ),
    .A3(_04509_),
    .A4(_04493_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09551_ (.A1(\delay_cycles[19] ),
    .A2(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09552_ (.I(\cycles_per_ms[19] ),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09553_ (.A1(_04507_),
    .A2(_04508_),
    .B1(_04511_),
    .B2(_04512_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09554_ (.I(\cycles_per_ms[17] ),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09555_ (.A1(_04509_),
    .A2(_04493_),
    .B(\delay_cycles[17] ),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09556_ (.A1(_04485_),
    .A2(_04494_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09557_ (.I(\cycles_per_ms[18] ),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09558_ (.A1(_04514_),
    .A2(_04495_),
    .A3(_04515_),
    .B1(_04516_),
    .B2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09559_ (.I(\cycles_per_ms[17] ),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09560_ (.A1(_04495_),
    .A2(_04515_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09561_ (.A1(_04509_),
    .A2(_04493_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09562_ (.I(\cycles_per_ms[16] ),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09563_ (.A1(_04519_),
    .A2(_04520_),
    .B1(_04521_),
    .B2(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09564_ (.I(\cycles_per_ms[19] ),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09565_ (.A1(\delay_cycles[19] ),
    .A2(_04510_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(_04522_),
    .A2(_04521_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09567_ (.A1(_04524_),
    .A2(_04525_),
    .B(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09568_ (.A1(_04513_),
    .A2(_04518_),
    .A3(_04523_),
    .A4(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09569_ (.I(\cycles_per_ms[15] ),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09570_ (.A1(_04487_),
    .A2(_04488_),
    .A3(_04492_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09571_ (.A1(\delay_cycles[15] ),
    .A2(_04530_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09572_ (.I(\delay_cycles[12] ),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09573_ (.I(_04491_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09574_ (.A1(_04532_),
    .A2(\delay_cycles[11] ),
    .A3(\delay_cycles[10] ),
    .A4(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09575_ (.A1(\delay_cycles[13] ),
    .A2(_04534_),
    .B(\delay_cycles[14] ),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09576_ (.A1(_04530_),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09577_ (.I(\cycles_per_ms[14] ),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09578_ (.I(_04537_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09579_ (.A1(_04529_),
    .A2(_04531_),
    .B1(_04536_),
    .B2(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09580_ (.I(\cycles_per_ms[15] ),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09581_ (.A1(_04486_),
    .A2(_04530_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09582_ (.I(\cycles_per_ms[13] ),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09583_ (.A1(_04488_),
    .A2(_04534_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09584_ (.I(\delay_cycles[11] ),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09585_ (.I(\delay_cycles[10] ),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09586_ (.A1(_04544_),
    .A2(_04545_),
    .A3(_04533_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09587_ (.A1(_04532_),
    .A2(_04546_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09588_ (.A1(_04542_),
    .A2(_04543_),
    .B1(_04547_),
    .B2(\cycles_per_ms[12] ),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09589_ (.A1(_04540_),
    .A2(_04541_),
    .B(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09590_ (.A1(\cycles_per_ms[14] ),
    .A2(_04530_),
    .A3(_04535_),
    .B1(_04543_),
    .B2(\cycles_per_ms[13] ),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09591_ (.I(\cycles_per_ms[12] ),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09592_ (.A1(_04551_),
    .A2(_04547_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09593_ (.A1(_04550_),
    .A2(_04552_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09594_ (.I(\cycles_per_ms[8] ),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09595_ (.I(\delay_cycles[8] ),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09596_ (.I(\delay_cycles[7] ),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_04556_),
    .A2(_04490_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09598_ (.A1(_04555_),
    .A2(_04557_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09599_ (.I(\cycles_per_ms[9] ),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09600_ (.A1(_04555_),
    .A2(_04556_),
    .A3(_04490_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09601_ (.A1(\delay_cycles[9] ),
    .A2(_04560_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09602_ (.A1(_04559_),
    .A2(_04561_),
    .B1(_04558_),
    .B2(\cycles_per_ms[8] ),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09603_ (.A1(_04545_),
    .A2(_04533_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09604_ (.A1(\cycles_per_ms[10] ),
    .A2(_04563_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09605_ (.I(\cycles_per_ms[10] ),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09606_ (.A1(_04565_),
    .A2(_04563_),
    .B1(_04561_),
    .B2(\cycles_per_ms[9] ),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09607_ (.A1(_04545_),
    .A2(_04533_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09608_ (.A1(_04544_),
    .A2(\cycles_per_ms[11] ),
    .A3(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09609_ (.A1(_04564_),
    .A2(_04566_),
    .A3(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09610_ (.A1(_04554_),
    .A2(_04558_),
    .B(_04562_),
    .C(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09611_ (.A1(_04539_),
    .A2(_04549_),
    .A3(_04553_),
    .A4(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09612_ (.I(\cycles_per_ms[7] ),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09613_ (.A1(_04556_),
    .A2(_04490_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09614_ (.I(\delay_cycles[4] ),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09615_ (.A1(\delay_cycles[5] ),
    .A2(_04574_),
    .A3(_04489_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09616_ (.A1(\delay_cycles[6] ),
    .A2(_04575_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09617_ (.I(\cycles_per_ms[6] ),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09618_ (.A1(_04572_),
    .A2(_04573_),
    .B1(_04576_),
    .B2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09619_ (.A1(_04574_),
    .A2(_04489_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09620_ (.A1(\delay_cycles[5] ),
    .A2(_04579_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09621_ (.A1(\cycles_per_ms[5] ),
    .A2(_04580_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09622_ (.A1(_04574_),
    .A2(_04489_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09623_ (.I(\delay_cycles[1] ),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09624_ (.I(\delay_cycles[0] ),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09625_ (.A1(\delay_cycles[2] ),
    .A2(_04583_),
    .A3(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09626_ (.A1(\delay_cycles[3] ),
    .A2(_04585_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09627_ (.I(\cycles_per_ms[3] ),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09628_ (.A1(\cycles_per_ms[4] ),
    .A2(_04582_),
    .B1(_04586_),
    .B2(_04587_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09629_ (.A1(_04583_),
    .A2(_04584_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09630_ (.A1(\delay_cycles[2] ),
    .A2(_04589_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09631_ (.A1(\cycles_per_ms[3] ),
    .A2(_04586_),
    .B1(_04590_),
    .B2(\cycles_per_ms[2] ),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09632_ (.I(\cycles_per_ms[5] ),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09633_ (.I(\cycles_per_ms[4] ),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09634_ (.A1(_04592_),
    .A2(_04580_),
    .B1(_04582_),
    .B2(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09635_ (.A1(_04588_),
    .A2(_04591_),
    .B(_04594_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09636_ (.A1(_04583_),
    .A2(_04584_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09637_ (.A1(\cycles_per_ms[1] ),
    .A2(_04596_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09638_ (.I(_04584_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09639_ (.A1(_04598_),
    .A2(\cycles_per_ms[0] ),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09640_ (.I(\cycles_per_ms[1] ),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09641_ (.A1(_04600_),
    .A2(_04596_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09642_ (.A1(_04597_),
    .A2(_04599_),
    .B(_04601_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09643_ (.I(\cycles_per_ms[2] ),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09644_ (.A1(_04603_),
    .A2(_04590_),
    .B(_04581_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09645_ (.A1(_04588_),
    .A2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09646_ (.A1(\cycles_per_ms[6] ),
    .A2(_04576_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09647_ (.A1(_04581_),
    .A2(_04595_),
    .B1(_04602_),
    .B2(_04605_),
    .C(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(_04572_),
    .A2(_04573_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09649_ (.A1(_04578_),
    .A2(_04607_),
    .B(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09650_ (.I(\cycles_per_ms[11] ),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09651_ (.A1(_04544_),
    .A2(_04567_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09652_ (.A1(_04610_),
    .A2(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09653_ (.A1(_04564_),
    .A2(_04566_),
    .A3(_04568_),
    .A4(_04562_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09654_ (.A1(_04610_),
    .A2(_04611_),
    .B(_04564_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09655_ (.A1(_04612_),
    .A2(_04613_),
    .A3(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09656_ (.A1(_04539_),
    .A2(_04549_),
    .A3(_04553_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(_04529_),
    .A2(_04531_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09658_ (.A1(_04550_),
    .A2(_04548_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09659_ (.A1(_04539_),
    .A2(_04618_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09660_ (.A1(_04571_),
    .A2(_04609_),
    .B1(_04615_),
    .B2(_04616_),
    .C1(_04617_),
    .C2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09661_ (.A1(_04507_),
    .A2(_04508_),
    .B1(_04520_),
    .B2(_04519_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09662_ (.A1(_04621_),
    .A2(_04523_),
    .B(_04513_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09663_ (.A1(_04524_),
    .A2(_04525_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09664_ (.A1(_04528_),
    .A2(_04620_),
    .B1(_04622_),
    .B2(_04623_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09665_ (.I(\cycles_per_ms[20] ),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09666_ (.A1(\delay_cycles[20] ),
    .A2(_04496_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09667_ (.A1(_04513_),
    .A2(_04518_),
    .A3(_04523_),
    .A4(_04527_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09668_ (.A1(_04597_),
    .A2(_04599_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09669_ (.I(\cycles_per_ms[0] ),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09670_ (.A1(_04598_),
    .A2(_04629_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09671_ (.A1(_04591_),
    .A2(_04601_),
    .A3(_04628_),
    .A4(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09672_ (.A1(_04606_),
    .A2(_04631_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09673_ (.A1(_04608_),
    .A2(_04594_),
    .A3(_04605_),
    .A4(_04632_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09674_ (.A1(_04578_),
    .A2(_04633_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09675_ (.A1(_04571_),
    .A2(_04634_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09676_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04627_),
    .B2(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09677_ (.A1(_04625_),
    .A2(_04626_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09678_ (.A1(_04505_),
    .A2(_04504_),
    .B1(_04624_),
    .B2(_04636_),
    .C(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09679_ (.A1(_04500_),
    .A2(_04501_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09680_ (.A1(_04484_),
    .A2(_04499_),
    .B1(_04506_),
    .B2(_04638_),
    .C(_04639_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09681_ (.A1(net142),
    .A2(_04252_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(_04250_),
    .A2(_04641_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09683_ (.A1(\delay_cycles[23] ),
    .A2(_04498_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09684_ (.A1(_04483_),
    .A2(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09685_ (.A1(\delay_cycles[23] ),
    .A2(_04498_),
    .B(_04642_),
    .C(_04644_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(_04253_),
    .A2(_04480_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09687_ (.A1(net143),
    .A2(_04641_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09688_ (.I(_04647_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09689_ (.I(_04648_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09690_ (.A1(\delay_counter[5] ),
    .A2(\delay_counter[4] ),
    .A3(\delay_counter[7] ),
    .A4(\delay_counter[6] ),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09691_ (.A1(\delay_counter[0] ),
    .A2(\delay_counter[1] ),
    .A3(\delay_counter[3] ),
    .A4(\delay_counter[2] ),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09692_ (.A1(_04650_),
    .A2(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09693_ (.A1(_01630_),
    .A2(_04258_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09694_ (.A1(_04254_),
    .A2(_04477_),
    .B1(_04649_),
    .B2(_04652_),
    .C(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_04646_),
    .A2(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09696_ (.A1(_04640_),
    .A2(_04645_),
    .B(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09697_ (.A1(_04469_),
    .A2(_04470_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09698_ (.A1(_04656_),
    .A2(_04657_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09699_ (.I(_04658_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09700_ (.A1(_04339_),
    .A2(_04473_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09701_ (.A1(_01769_),
    .A2(_04325_),
    .A3(_01896_),
    .A4(_01988_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09702_ (.A1(_01800_),
    .A2(_01833_),
    .B1(_01960_),
    .B2(_04444_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09703_ (.A1(_01800_),
    .A2(_01833_),
    .B1(_01959_),
    .B2(_04444_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09704_ (.I(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09705_ (.A1(_04661_),
    .A2(_04662_),
    .A3(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09706_ (.A1(_04250_),
    .A2(_04251_),
    .A3(_04256_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09707_ (.A1(_04478_),
    .A2(_04666_),
    .A3(_04649_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09708_ (.A1(_04322_),
    .A2(_04333_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09709_ (.A1(_04353_),
    .A2(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09710_ (.A1(_04276_),
    .A2(_04297_),
    .A3(_04311_),
    .A4(_04344_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09711_ (.A1(_04276_),
    .A2(_04297_),
    .A3(_04311_),
    .A4(_04344_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09712_ (.A1(_04670_),
    .A2(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09713_ (.A1(_04286_),
    .A2(_04667_),
    .A3(_04669_),
    .A4(_04672_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09714_ (.I(_04648_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09715_ (.A1(_04480_),
    .A2(_04674_),
    .B(single_step),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09716_ (.A1(_04412_),
    .A2(_01240_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09717_ (.I(single_step),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09718_ (.A1(_04677_),
    .A2(_01244_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09719_ (.A1(_04413_),
    .A2(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09720_ (.A1(_04673_),
    .A2(_04675_),
    .A3(_04676_),
    .A4(_04679_),
    .Z(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09721_ (.A1(_04660_),
    .A2(_04665_),
    .B1(_04680_),
    .B2(_04388_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09722_ (.A1(_04659_),
    .A2(_04681_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09723_ (.A1(_04256_),
    .A2(_04659_),
    .B(_04682_),
    .C(_02010_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09724_ (.A1(_04251_),
    .A2(_04659_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09725_ (.A1(_04388_),
    .A2(_04473_),
    .A3(_04665_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09726_ (.I(_04250_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09727_ (.A1(_04685_),
    .A2(_04257_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09728_ (.A1(_04686_),
    .A2(_04676_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09729_ (.A1(_04667_),
    .A2(_04687_),
    .B(_04673_),
    .C(_04324_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09730_ (.A1(_04658_),
    .A2(_04684_),
    .A3(_04688_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09731_ (.A1(_03594_),
    .A2(_04683_),
    .A3(_04689_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09732_ (.A1(_01624_),
    .A2(_01590_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09733_ (.A1(_01189_),
    .A2(_01194_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09734_ (.A1(\cycles_per_ms[19] ),
    .A2(_04517_),
    .A3(_04514_),
    .A4(\cycles_per_ms[16] ),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09735_ (.A1(\cycles_per_ms[23] ),
    .A2(\cycles_per_ms[22] ),
    .A3(\cycles_per_ms[21] ),
    .A4(\cycles_per_ms[20] ),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09736_ (.A1(_04692_),
    .A2(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09737_ (.A1(\cycles_per_ms[11] ),
    .A2(_04565_),
    .A3(_04559_),
    .A4(_04554_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09738_ (.A1(_04540_),
    .A2(_04537_),
    .A3(_04542_),
    .A4(_04551_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09739_ (.A1(_04587_),
    .A2(_04603_),
    .A3(_04600_),
    .A4(_04629_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09740_ (.A1(\cycles_per_ms[7] ),
    .A2(_04577_),
    .A3(_04592_),
    .A4(_04593_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09741_ (.A1(_04695_),
    .A2(_04696_),
    .A3(_04697_),
    .A4(_04698_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09742_ (.A1(_01168_),
    .A2(_01969_),
    .B1(_04694_),
    .B2(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09743_ (.A1(_04691_),
    .A2(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09744_ (.A1(_04678_),
    .A2(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09745_ (.A1(_04690_),
    .A2(_04702_),
    .B(_04675_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09746_ (.A1(_04403_),
    .A2(_04656_),
    .A3(_04703_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09747_ (.A1(_04685_),
    .A2(_04659_),
    .B(_04704_),
    .C(_02010_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09748_ (.A1(_03625_),
    .A2(_01241_),
    .B(\intr[0] ),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09749_ (.A1(_03619_),
    .A2(_04277_),
    .B(_04705_),
    .C(_04467_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09750_ (.A1(_03618_),
    .A2(_04361_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09751_ (.A1(\intr_enable[0] ),
    .A2(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09752_ (.I(_04336_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09753_ (.A1(_01727_),
    .A2(_04706_),
    .B(_04707_),
    .C(_04708_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09754_ (.A1(\intr_enable[1] ),
    .A2(_04706_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09755_ (.A1(_03623_),
    .A2(_04706_),
    .B(_04709_),
    .C(_04708_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09756_ (.A1(edge_interrupts),
    .A2(_04474_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09757_ (.A1(_04312_),
    .A2(_04475_),
    .B(_04710_),
    .C(_04708_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09758_ (.A1(_01644_),
    .A2(_04387_),
    .A3(_04254_),
    .A4(_04686_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09759_ (.I(_04711_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09760_ (.I0(\exec.memory_input[0] ),
    .I1(_04276_),
    .S(_04712_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09761_ (.I(_04713_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09762_ (.I0(\exec.memory_input[1] ),
    .I1(_04286_),
    .S(_04712_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09763_ (.I(_04714_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09764_ (.I(_04711_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09765_ (.I0(\exec.memory_input[2] ),
    .I1(_04297_),
    .S(_04715_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09766_ (.I(_04716_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09767_ (.I0(\exec.memory_input[3] ),
    .I1(_04311_),
    .S(_04715_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09768_ (.I(_04717_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09769_ (.I0(\exec.memory_input[4] ),
    .I1(_04322_),
    .S(_04715_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09770_ (.I(_04718_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09771_ (.I0(\exec.memory_input[5] ),
    .I1(_04333_),
    .S(_04715_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09772_ (.I(_04719_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09773_ (.A1(\exec.memory_input[6] ),
    .A2(_04712_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09774_ (.A1(_04344_),
    .A2(_04712_),
    .B(_04720_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09775_ (.I0(\exec.memory_input[7] ),
    .I1(_04353_),
    .S(_04711_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09776_ (.I(_04721_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09777_ (.A1(single_step),
    .A2(_04262_),
    .A3(_04474_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09778_ (.A1(_03623_),
    .A2(_04475_),
    .B(_04722_),
    .C(_04708_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09779_ (.A1(_04468_),
    .A2(_01179_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09780_ (.A1(_04412_),
    .A2(_04477_),
    .B(_03620_),
    .C(_02127_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09781_ (.I(_04723_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09782_ (.A1(_01224_),
    .A2(_01245_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09783_ (.A1(_04413_),
    .A2(_01238_),
    .B1(_04725_),
    .B2(_04666_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09784_ (.A1(_00764_),
    .A2(_04724_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09785_ (.A1(_04724_),
    .A2(_04726_),
    .B(_04727_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09786_ (.I(_04724_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09787_ (.A1(_04412_),
    .A2(_04666_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09788_ (.I(_04729_),
    .Z(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09789_ (.I(_04723_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09790_ (.I(_04729_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09791_ (.A1(_03889_),
    .A2(_04732_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09792_ (.A1(net128),
    .A2(_04730_),
    .B(_04731_),
    .C(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09793_ (.A1(_00757_),
    .A2(_04728_),
    .B(_04734_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09794_ (.A1(_01762_),
    .A2(_04732_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09795_ (.A1(_04376_),
    .A2(_04730_),
    .B(_04731_),
    .C(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09796_ (.A1(_00756_),
    .A2(_04728_),
    .B(_04736_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09797_ (.A1(_01795_),
    .A2(_04732_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09798_ (.A1(net257),
    .A2(_04730_),
    .B(_04731_),
    .C(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09799_ (.A1(_03098_),
    .A2(_04728_),
    .B(_04738_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09800_ (.I(_04729_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09801_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09802_ (.I(_04723_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09803_ (.A1(_01827_),
    .A2(_04732_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09804_ (.A1(net153),
    .A2(_04740_),
    .B(_04741_),
    .C(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09805_ (.A1(_02813_),
    .A2(_04728_),
    .B(_04743_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09806_ (.I(_04731_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09807_ (.A1(_01859_),
    .A2(_04739_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09808_ (.A1(_04406_),
    .A2(_04740_),
    .B(_04741_),
    .C(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09809_ (.A1(_02760_),
    .A2(_04744_),
    .B(_04746_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09810_ (.A1(_01891_),
    .A2(_04739_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09811_ (.A1(_04417_),
    .A2(_04740_),
    .B(_04741_),
    .C(_04747_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09812_ (.A1(_01173_),
    .A2(_04744_),
    .B(_04748_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09813_ (.I(net189),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09814_ (.A1(_04413_),
    .A2(_04666_),
    .B(_01125_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09815_ (.A1(_04423_),
    .A2(_04730_),
    .B(_04724_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09816_ (.A1(_04749_),
    .A2(_04744_),
    .B1(_04750_),
    .B2(_04751_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09817_ (.I(net190),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09818_ (.A1(_03737_),
    .A2(_04739_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09819_ (.A1(net157),
    .A2(_04740_),
    .B(_04741_),
    .C(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09820_ (.A1(_04752_),
    .A2(_04744_),
    .B(_04754_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09821_ (.A1(net232),
    .A2(_02033_),
    .A3(_04481_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09822_ (.A1(_04375_),
    .A2(_04440_),
    .A3(_04646_),
    .B(_04755_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09823_ (.A1(_01694_),
    .A2(_04362_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09824_ (.I(_04756_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09825_ (.I(_04757_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09826_ (.I(_04757_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09827_ (.A1(_04629_),
    .A2(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09828_ (.I(_04336_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09829_ (.A1(_01727_),
    .A2(_04758_),
    .B(_04760_),
    .C(_04761_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09830_ (.I(_04756_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09831_ (.A1(_04600_),
    .A2(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09832_ (.A1(_03623_),
    .A2(_04758_),
    .B(_04763_),
    .C(_04761_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09833_ (.A1(_04603_),
    .A2(_04762_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09834_ (.A1(_04299_),
    .A2(_04758_),
    .B(_04764_),
    .C(_04761_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09835_ (.A1(_04587_),
    .A2(_04762_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09836_ (.A1(_04312_),
    .A2(_04758_),
    .B(_04765_),
    .C(_04761_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09837_ (.A1(_01694_),
    .A2(_04362_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09838_ (.I(_04766_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09839_ (.I(_04766_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09840_ (.I(_04768_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09841_ (.A1(_04593_),
    .A2(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09842_ (.A1(_04325_),
    .A2(_04767_),
    .B(_04770_),
    .C(_02010_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09843_ (.A1(_04592_),
    .A2(_04762_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09844_ (.A1(_01896_),
    .A2(_04759_),
    .B(_04771_),
    .C(_03569_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09845_ (.A1(_04577_),
    .A2(_04757_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09846_ (.A1(_01960_),
    .A2(_04759_),
    .B(_04772_),
    .C(_03569_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09847_ (.A1(_04572_),
    .A2(_04757_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09848_ (.A1(_04356_),
    .A2(_04759_),
    .B(_04773_),
    .C(_03569_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09849_ (.A1(_04354_),
    .A2(_04766_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09850_ (.I(_04774_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09851_ (.I(_04374_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09852_ (.A1(_04554_),
    .A2(_04767_),
    .B1(_04775_),
    .B2(net65),
    .C(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09853_ (.I(_04777_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09854_ (.A1(_04559_),
    .A2(_04767_),
    .B1(_04775_),
    .B2(net66),
    .C(_03262_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09855_ (.I(_04778_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09856_ (.A1(_04565_),
    .A2(_04767_),
    .B1(_04775_),
    .B2(net44),
    .C(_03262_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09857_ (.I(_04779_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09858_ (.I(_04774_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09859_ (.A1(_04610_),
    .A2(_04769_),
    .B1(_04780_),
    .B2(net45),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09860_ (.A1(_04468_),
    .A2(_04781_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09861_ (.A1(_04551_),
    .A2(_04769_),
    .B1(_04780_),
    .B2(net46),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09862_ (.A1(_04468_),
    .A2(_04782_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09863_ (.A1(_04542_),
    .A2(_04769_),
    .B1(_04775_),
    .B2(net47),
    .C(_03262_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09864_ (.I(_04783_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09865_ (.I(_03281_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09866_ (.I(_04768_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09867_ (.A1(_04537_),
    .A2(_04785_),
    .B1(_04780_),
    .B2(net48),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09868_ (.A1(_04784_),
    .A2(_04786_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09869_ (.A1(_04540_),
    .A2(_04785_),
    .B1(_04780_),
    .B2(net49),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09870_ (.A1(_04784_),
    .A2(_04787_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09871_ (.I(_04774_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09872_ (.A1(\cycles_per_ms[16] ),
    .A2(_04785_),
    .B1(_04788_),
    .B2(net50),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09873_ (.A1(_04784_),
    .A2(_04789_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09874_ (.A1(_04514_),
    .A2(_04785_),
    .B1(_04788_),
    .B2(net51),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09875_ (.A1(_04784_),
    .A2(_04790_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09876_ (.I(_03281_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09877_ (.I(_04766_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09878_ (.A1(_04517_),
    .A2(_04792_),
    .B1(_04788_),
    .B2(net52),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09879_ (.A1(_04791_),
    .A2(_04793_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09880_ (.A1(_04524_),
    .A2(_04792_),
    .B1(_04788_),
    .B2(net53),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09881_ (.A1(_04791_),
    .A2(_04794_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09882_ (.I(_04774_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09883_ (.A1(\cycles_per_ms[20] ),
    .A2(_04792_),
    .B1(_04795_),
    .B2(net55),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09884_ (.A1(_04791_),
    .A2(_04796_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09885_ (.A1(_04505_),
    .A2(_04792_),
    .B1(_04795_),
    .B2(net56),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09886_ (.A1(_04791_),
    .A2(_04797_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09887_ (.I(_03261_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09888_ (.I(_04798_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09889_ (.A1(_04500_),
    .A2(_04768_),
    .B1(_04795_),
    .B2(net57),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09890_ (.A1(_04799_),
    .A2(_04800_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09891_ (.A1(_04483_),
    .A2(_04768_),
    .B1(_04795_),
    .B2(net58),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09892_ (.A1(_04799_),
    .A2(_04801_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09893_ (.I(_04678_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09894_ (.A1(_04802_),
    .A2(_04701_),
    .B(_04690_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09895_ (.A1(_01624_),
    .A2(_01590_),
    .B(_04648_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _09896_ (.A1(_04338_),
    .A2(_04803_),
    .A3(_04804_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09897_ (.I(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09898_ (.A1(_04640_),
    .A2(_04645_),
    .A3(_04806_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09899_ (.I(_04807_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09900_ (.A1(_04598_),
    .A2(_04808_),
    .B(_03183_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09901_ (.A1(_04598_),
    .A2(_04806_),
    .B(_04809_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09902_ (.I(_04805_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09903_ (.I(_04810_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09904_ (.I(_04596_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09905_ (.A1(_04583_),
    .A2(_04811_),
    .B1(_04808_),
    .B2(_04812_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09906_ (.A1(_04799_),
    .A2(_04813_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09907_ (.I(_04590_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09908_ (.A1(\delay_cycles[2] ),
    .A2(_04811_),
    .B1(_04808_),
    .B2(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09909_ (.A1(_04799_),
    .A2(_04815_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09910_ (.I(_04798_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09911_ (.I(_04586_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09912_ (.A1(\delay_cycles[3] ),
    .A2(_04811_),
    .B1(_04808_),
    .B2(_04817_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09913_ (.A1(_04816_),
    .A2(_04818_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09914_ (.I(_04807_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09915_ (.I(_04819_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09916_ (.I(_04582_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09917_ (.A1(_04574_),
    .A2(_04811_),
    .B1(_04820_),
    .B2(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09918_ (.A1(_04816_),
    .A2(_04822_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09919_ (.I(_04805_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09920_ (.I(_04823_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09921_ (.I(_04580_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09922_ (.A1(\delay_cycles[5] ),
    .A2(_04824_),
    .B1(_04820_),
    .B2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09923_ (.A1(_04816_),
    .A2(_04826_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09924_ (.I(_04576_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09925_ (.A1(\delay_cycles[6] ),
    .A2(_04824_),
    .B1(_04820_),
    .B2(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09926_ (.A1(_04816_),
    .A2(_04828_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09927_ (.I(_04798_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09928_ (.I(_04573_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09929_ (.A1(_04556_),
    .A2(_04824_),
    .B1(_04820_),
    .B2(_04830_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09930_ (.A1(_04829_),
    .A2(_04831_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09931_ (.I(_04819_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09932_ (.A1(_04555_),
    .A2(_04557_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09933_ (.A1(_04555_),
    .A2(_04824_),
    .B1(_04832_),
    .B2(_04833_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09934_ (.A1(_04829_),
    .A2(_04834_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09935_ (.I(_04823_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09936_ (.A1(\delay_cycles[9] ),
    .A2(_04560_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09937_ (.A1(\delay_cycles[9] ),
    .A2(_04835_),
    .B1(_04832_),
    .B2(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09938_ (.A1(_04829_),
    .A2(_04837_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09939_ (.I(_04563_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09940_ (.A1(_04545_),
    .A2(_04835_),
    .B1(_04832_),
    .B2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09941_ (.A1(_04829_),
    .A2(_04839_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09942_ (.I(_04798_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09943_ (.I(_04611_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09944_ (.A1(_04544_),
    .A2(_04835_),
    .B1(_04832_),
    .B2(_04841_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09945_ (.A1(_04840_),
    .A2(_04842_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09946_ (.I(_04819_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09947_ (.A1(_04532_),
    .A2(_04546_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09948_ (.A1(_04532_),
    .A2(_04835_),
    .B1(_04843_),
    .B2(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09949_ (.A1(_04840_),
    .A2(_04845_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09950_ (.I(_04823_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09951_ (.A1(\delay_cycles[13] ),
    .A2(_04534_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09952_ (.A1(\delay_cycles[13] ),
    .A2(_04846_),
    .B1(_04843_),
    .B2(_04847_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09953_ (.A1(_04840_),
    .A2(_04848_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09954_ (.A1(\delay_cycles[14] ),
    .A2(_04846_),
    .B1(_04843_),
    .B2(_04536_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09955_ (.A1(_04840_),
    .A2(_04849_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09956_ (.I(_02004_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09957_ (.A1(\delay_cycles[15] ),
    .A2(_04846_),
    .B1(_04843_),
    .B2(_04531_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09958_ (.A1(_04850_),
    .A2(_04851_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09959_ (.I(_04819_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09960_ (.A1(_04509_),
    .A2(_04846_),
    .B1(_04852_),
    .B2(_04521_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09961_ (.A1(_04850_),
    .A2(_04853_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09962_ (.I(_04823_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09963_ (.A1(\delay_cycles[17] ),
    .A2(_04854_),
    .B1(_04852_),
    .B2(_04520_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09964_ (.A1(_04850_),
    .A2(_04855_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09965_ (.A1(_04485_),
    .A2(_04854_),
    .B1(_04852_),
    .B2(_04508_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09966_ (.A1(_04850_),
    .A2(_04856_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09967_ (.I(_02004_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09968_ (.A1(\delay_cycles[19] ),
    .A2(_04854_),
    .B1(_04852_),
    .B2(_04511_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09969_ (.A1(_04857_),
    .A2(_04858_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09970_ (.I(_04807_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09971_ (.A1(\delay_cycles[20] ),
    .A2(_04854_),
    .B1(_04859_),
    .B2(_04626_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09972_ (.A1(_04857_),
    .A2(_04860_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09973_ (.A1(\delay_cycles[21] ),
    .A2(_04810_),
    .B1(_04859_),
    .B2(_04503_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09974_ (.A1(_04857_),
    .A2(_04861_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09975_ (.I(_04501_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09976_ (.A1(\delay_cycles[22] ),
    .A2(_04810_),
    .B1(_04859_),
    .B2(_04862_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09977_ (.A1(_04857_),
    .A2(_04863_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09978_ (.A1(\delay_cycles[23] ),
    .A2(_04810_),
    .B1(_04859_),
    .B2(_04499_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09979_ (.A1(_03627_),
    .A2(_04864_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09980_ (.I(_01633_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09981_ (.I(_04865_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09982_ (.I(_04865_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_02031_),
    .A2(_04867_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09984_ (.A1(_04866_),
    .A2(_01738_),
    .B(_04868_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09985_ (.I(_04865_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09986_ (.I(_04865_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09987_ (.A1(_04870_),
    .A2(_01782_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09988_ (.A1(_02994_),
    .A2(_04869_),
    .B(_04871_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09989_ (.A1(_02041_),
    .A2(_04867_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09990_ (.A1(_04866_),
    .A2(_01837_),
    .B(_04872_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09991_ (.A1(_04870_),
    .A2(_01835_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09992_ (.A1(_02998_),
    .A2(_04869_),
    .B(_04873_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09993_ (.A1(_02051_),
    .A2(_04867_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09994_ (.A1(_04866_),
    .A2(_01878_),
    .B(_04874_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09995_ (.A1(_02056_),
    .A2(_04867_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09996_ (.A1(_04866_),
    .A2(_01904_),
    .B(_04875_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09997_ (.A1(_04870_),
    .A2(_01949_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09998_ (.A1(_03007_),
    .A2(_04869_),
    .B(_04876_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09999_ (.A1(_04870_),
    .A2(_01968_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10000_ (.A1(_03009_),
    .A2(_04869_),
    .B(_04877_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10001_ (.A1(wb_write_ack),
    .A2(_04354_),
    .B(_01628_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10002_ (.A1(_03627_),
    .A2(_04878_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10003_ (.A1(_04691_),
    .A2(_04647_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10004_ (.A1(\delay_counter[0] ),
    .A2(_04647_),
    .B1(_04879_),
    .B2(_00841_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10005_ (.A1(_04640_),
    .A2(_04645_),
    .B(_04805_),
    .C(_01644_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10006_ (.I(_04881_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10007_ (.I0(\delay_counter[0] ),
    .I1(_04880_),
    .S(_04882_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10008_ (.I(_04883_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10009_ (.I(_04881_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10010_ (.I(_04879_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10011_ (.A1(\delay_counter[1] ),
    .A2(_04647_),
    .B1(_04885_),
    .B2(_00876_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10012_ (.A1(_04880_),
    .A2(_04886_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10013_ (.I(_04881_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10014_ (.A1(\delay_counter[1] ),
    .A2(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10015_ (.A1(_04884_),
    .A2(_04887_),
    .B(_04889_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10016_ (.A1(_04880_),
    .A2(_04886_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10017_ (.A1(\delay_counter[2] ),
    .A2(_04648_),
    .B1(_04885_),
    .B2(_00919_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10018_ (.A1(_04890_),
    .A2(_04891_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10019_ (.A1(\delay_counter[2] ),
    .A2(_04888_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10020_ (.A1(_04884_),
    .A2(_04892_),
    .B(_04893_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10021_ (.A1(_04890_),
    .A2(_04891_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10022_ (.A1(\delay_counter[3] ),
    .A2(_04649_),
    .B1(_04885_),
    .B2(_00983_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10023_ (.A1(_04894_),
    .A2(_04895_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10024_ (.A1(\delay_counter[3] ),
    .A2(_04888_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10025_ (.A1(_04884_),
    .A2(_04896_),
    .B(_04897_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10026_ (.A1(_04894_),
    .A2(_04895_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10027_ (.I(_04885_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10028_ (.A1(\delay_counter[4] ),
    .A2(_04649_),
    .B1(_04899_),
    .B2(_01027_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10029_ (.A1(_04898_),
    .A2(_04900_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10030_ (.I0(\delay_counter[4] ),
    .I1(_04901_),
    .S(_04882_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10031_ (.I(_04902_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10032_ (.A1(_04894_),
    .A2(_04895_),
    .A3(_04900_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10033_ (.A1(\delay_counter[5] ),
    .A2(_04674_),
    .B1(_04899_),
    .B2(_01075_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10034_ (.A1(_04903_),
    .A2(_04904_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10035_ (.A1(\delay_counter[5] ),
    .A2(_04882_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10036_ (.A1(_04884_),
    .A2(_04905_),
    .B(_04906_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10037_ (.A1(_04903_),
    .A2(_04904_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10038_ (.A1(\delay_counter[6] ),
    .A2(_04674_),
    .B1(_04899_),
    .B2(_01123_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10039_ (.A1(_04907_),
    .A2(_04908_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10040_ (.I0(\delay_counter[6] ),
    .I1(_04909_),
    .S(_04881_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10041_ (.I(_04910_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10042_ (.A1(_04903_),
    .A2(_04904_),
    .A3(_04908_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10043_ (.A1(\delay_counter[7] ),
    .A2(_04674_),
    .B1(_04899_),
    .B2(_01169_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10044_ (.A1(_04911_),
    .A2(_04912_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10045_ (.A1(\delay_counter[7] ),
    .A2(_04882_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10046_ (.A1(_04888_),
    .A2(_04913_),
    .B(_04914_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10047_ (.I(_00842_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10048_ (.A1(net38),
    .A2(net39),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10049_ (.A1(net22),
    .A2(net21),
    .A3(net24),
    .A4(net23),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10050_ (.A1(net41),
    .A2(net40),
    .A3(net20),
    .A4(net19),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10051_ (.A1(_04917_),
    .A2(_04918_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10052_ (.A1(net37),
    .A2(_04919_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10053_ (.A1(net36),
    .A2(_04916_),
    .A3(_04920_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10054_ (.I(net35),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10055_ (.A1(net31),
    .A2(net30),
    .A3(net33),
    .A4(net32),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10056_ (.A1(net26),
    .A2(net25),
    .A3(net28),
    .A4(net27),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10057_ (.A1(net34),
    .A2(_01655_),
    .A3(_04923_),
    .A4(_04924_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10058_ (.A1(_04922_),
    .A2(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10059_ (.A1(_04921_),
    .A2(_04926_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10060_ (.I(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10061_ (.A1(net18),
    .A2(net29),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10062_ (.A1(_04923_),
    .A2(_04924_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10063_ (.A1(net36),
    .A2(net38),
    .A3(net39),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10064_ (.A1(_04931_),
    .A2(_04920_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(_04922_),
    .A2(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10066_ (.A1(net34),
    .A2(_04929_),
    .A3(_04930_),
    .A4(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10067_ (.I(_04934_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10068_ (.A1(net34),
    .A2(_04922_),
    .A3(_04929_),
    .A4(_04930_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10069_ (.I(_04932_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10070_ (.A1(_04936_),
    .A2(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10071_ (.I(_04938_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10072_ (.A1(_01197_),
    .A2(_04935_),
    .B1(_04939_),
    .B2(net128),
    .C(_04139_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10073_ (.A1(_04933_),
    .A2(_04925_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10074_ (.A1(_04258_),
    .A2(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10075_ (.A1(_04932_),
    .A2(_04926_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10076_ (.I(_04943_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10077_ (.A1(net37),
    .A2(_04917_),
    .A3(_04918_),
    .A4(_04931_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10078_ (.A1(_04922_),
    .A2(_04925_),
    .A3(_04945_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10079_ (.A1(_01700_),
    .A2(_04944_),
    .B1(_04946_),
    .B2(\intr[0] ),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10080_ (.I(_04921_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10081_ (.A1(_04936_),
    .A2(_04948_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10082_ (.I(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10083_ (.A1(_04936_),
    .A2(_04945_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10084_ (.A1(_04629_),
    .A2(_04950_),
    .B1(_04951_),
    .B2(\intr_enable[0] ),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10085_ (.A1(_04940_),
    .A2(_04942_),
    .A3(_04947_),
    .A4(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10086_ (.A1(_04915_),
    .A2(_04928_),
    .B(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10087_ (.A1(net68),
    .A2(_01627_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10088_ (.I(_04955_),
    .Z(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10089_ (.I(_04956_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10090_ (.A1(net161),
    .A2(_04957_),
    .B(_04429_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10091_ (.A1(_04954_),
    .A2(_04958_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10092_ (.A1(_01211_),
    .A2(_04935_),
    .B1(_04951_),
    .B2(\intr_enable[1] ),
    .C(_04139_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(single_step),
    .A2(_04941_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10094_ (.I(_04938_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10095_ (.A1(_04376_),
    .A2(_04961_),
    .B1(_04944_),
    .B2(_01114_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10096_ (.I(_04949_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10097_ (.A1(_04600_),
    .A2(_04963_),
    .B1(_04946_),
    .B2(\intr[1] ),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10098_ (.A1(_04959_),
    .A2(_04960_),
    .A3(_04962_),
    .A4(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10099_ (.A1(_00877_),
    .A2(_04928_),
    .B(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10100_ (.A1(net172),
    .A2(_04957_),
    .B(_04429_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10101_ (.A1(_04966_),
    .A2(_04967_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10102_ (.I(net177),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10103_ (.I(_04934_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10104_ (.A1(_04603_),
    .A2(_04963_),
    .B1(_04944_),
    .B2(_01133_),
    .C1(net257),
    .C2(_04939_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10105_ (.A1(_04956_),
    .A2(_04970_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10106_ (.A1(_01228_),
    .A2(_04969_),
    .B1(_04941_),
    .B2(_04281_),
    .C(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10107_ (.I(_04927_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_04100_),
    .A2(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10109_ (.A1(_04968_),
    .A2(_04141_),
    .B1(_04972_),
    .B2(_04974_),
    .C(_04776_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10110_ (.I(net178),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10111_ (.I(_04955_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10112_ (.A1(_04587_),
    .A2(_04963_),
    .B1(_04943_),
    .B2(_01255_),
    .C1(net153),
    .C2(_04939_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10113_ (.A1(_04976_),
    .A2(_04977_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10114_ (.A1(_01191_),
    .A2(_04935_),
    .B1(_04941_),
    .B2(edge_interrupts),
    .C(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(_04103_),
    .A2(_04973_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10116_ (.A1(_04975_),
    .A2(_04141_),
    .B1(_04979_),
    .B2(_04980_),
    .C(_04776_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10117_ (.A1(_01215_),
    .A2(_04935_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10118_ (.A1(_04593_),
    .A2(_04963_),
    .B1(_04944_),
    .B2(_00778_),
    .C1(_04406_),
    .C2(_04939_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10119_ (.A1(_04956_),
    .A2(_04981_),
    .A3(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10120_ (.A1(_01027_),
    .A2(_04928_),
    .B(_04983_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10121_ (.A1(net179),
    .A2(_04957_),
    .B(_04429_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10122_ (.A1(_04984_),
    .A2(_04985_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10123_ (.I(_04949_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10124_ (.A1(_04417_),
    .A2(_04961_),
    .B1(_04986_),
    .B2(_04592_),
    .C(_04140_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10125_ (.A1(_01233_),
    .A2(_04969_),
    .B1(_04928_),
    .B2(_01075_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10126_ (.A1(net180),
    .A2(_04957_),
    .B(_03183_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10127_ (.A1(_04987_),
    .A2(_04988_),
    .B(_04989_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10128_ (.I(net181),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10129_ (.A1(_04423_),
    .A2(_04961_),
    .B1(_04986_),
    .B2(_04577_),
    .C(_04140_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10130_ (.A1(_01217_),
    .A2(_04969_),
    .B1(_04973_),
    .B2(_01125_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10131_ (.A1(_04990_),
    .A2(_04141_),
    .B1(_04991_),
    .B2(_04992_),
    .C(_04776_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10132_ (.A1(net157),
    .A2(_04961_),
    .B1(_04986_),
    .B2(_04572_),
    .C(_04140_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10133_ (.I(_01169_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10134_ (.A1(_01216_),
    .A2(_04969_),
    .B1(_04973_),
    .B2(_04994_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10135_ (.I(_04955_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10136_ (.A1(net182),
    .A2(_04996_),
    .B(_03183_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10137_ (.A1(_04993_),
    .A2(_04995_),
    .B(_04997_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10138_ (.I(_04139_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10139_ (.I(_04998_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10140_ (.A1(net183),
    .A2(_04999_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10141_ (.I(_04986_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10142_ (.A1(_04554_),
    .A2(_04996_),
    .A3(_05001_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10143_ (.A1(_05000_),
    .A2(_05002_),
    .B(_04472_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10144_ (.A1(net184),
    .A2(_04999_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10145_ (.A1(_04559_),
    .A2(_04996_),
    .A3(_05001_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10146_ (.A1(_05003_),
    .A2(_05004_),
    .B(_04472_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10147_ (.A1(net162),
    .A2(_04999_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10148_ (.A1(_04565_),
    .A2(_04996_),
    .A3(_05001_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10149_ (.A1(_05005_),
    .A2(_05006_),
    .B(_04472_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10150_ (.A1(net163),
    .A2(_04999_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10151_ (.I(_04976_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10152_ (.A1(_04610_),
    .A2(_05008_),
    .A3(_05001_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10153_ (.I(_04288_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10154_ (.A1(_05007_),
    .A2(_05009_),
    .B(_05010_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10155_ (.I(_04998_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10156_ (.A1(net164),
    .A2(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10157_ (.I(_04950_),
    .Z(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10158_ (.A1(_04551_),
    .A2(_05008_),
    .A3(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10159_ (.A1(_05012_),
    .A2(_05014_),
    .B(_05010_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10160_ (.A1(net165),
    .A2(_05011_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10161_ (.A1(_04542_),
    .A2(_05008_),
    .A3(_05013_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10162_ (.A1(_05015_),
    .A2(_05016_),
    .B(_05010_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10163_ (.A1(net166),
    .A2(_05011_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10164_ (.A1(_04537_),
    .A2(_05008_),
    .A3(_05013_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10165_ (.A1(_05017_),
    .A2(_05018_),
    .B(_05010_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10166_ (.A1(net167),
    .A2(_05011_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10167_ (.I(_04976_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10168_ (.A1(_04540_),
    .A2(_05020_),
    .A3(_05013_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10169_ (.I(_04288_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10170_ (.A1(_05019_),
    .A2(_05021_),
    .B(_05022_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10171_ (.I(_04998_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10172_ (.A1(net168),
    .A2(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10173_ (.I(_04950_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10174_ (.A1(\cycles_per_ms[16] ),
    .A2(_05020_),
    .A3(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10175_ (.A1(_05024_),
    .A2(_05026_),
    .B(_05022_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10176_ (.A1(net169),
    .A2(_05023_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10177_ (.A1(_04514_),
    .A2(_05020_),
    .A3(_05025_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10178_ (.A1(_05027_),
    .A2(_05028_),
    .B(_05022_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10179_ (.A1(net170),
    .A2(_05023_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10180_ (.A1(_04517_),
    .A2(_05020_),
    .A3(_05025_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10181_ (.A1(_05029_),
    .A2(_05030_),
    .B(_05022_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10182_ (.A1(net171),
    .A2(_05023_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10183_ (.I(_04976_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10184_ (.A1(_04524_),
    .A2(_05032_),
    .A3(_05025_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10185_ (.I(_04288_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10186_ (.A1(_05031_),
    .A2(_05033_),
    .B(_05034_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10187_ (.I(_04998_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10188_ (.A1(net173),
    .A2(_05035_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10189_ (.I(_04950_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10190_ (.A1(\cycles_per_ms[20] ),
    .A2(_05032_),
    .A3(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10191_ (.A1(_05036_),
    .A2(_05038_),
    .B(_05034_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10192_ (.A1(net174),
    .A2(_05035_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10193_ (.A1(_04505_),
    .A2(_05032_),
    .A3(_05037_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10194_ (.A1(_05039_),
    .A2(_05040_),
    .B(_05034_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10195_ (.A1(net175),
    .A2(_05035_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10196_ (.A1(_04500_),
    .A2(_05032_),
    .A3(_05037_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10197_ (.A1(_05041_),
    .A2(_05042_),
    .B(_05034_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(net176),
    .A2(_05035_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10199_ (.A1(_04483_),
    .A2(_04956_),
    .A3(_05037_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10200_ (.A1(_05043_),
    .A2(_05044_),
    .B(_02005_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10201_ (.A1(_03635_),
    .A2(_03701_),
    .A3(_03994_),
    .A4(_03192_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10202_ (.A1(_03202_),
    .A2(_03990_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10203_ (.A1(_04185_),
    .A2(_05045_),
    .A3(_05046_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10204_ (.I(_05047_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10205_ (.A1(\stack[12][0] ),
    .A2(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10206_ (.I(_05045_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10207_ (.I(_05046_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10208_ (.A1(_04191_),
    .A2(_05050_),
    .B1(_05051_),
    .B2(_04167_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10209_ (.A1(_05049_),
    .A2(_05052_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10210_ (.I(_03868_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10211_ (.I(_05051_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10212_ (.I(_05054_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10213_ (.A1(_04218_),
    .A2(_05050_),
    .B1(_05048_),
    .B2(\stack[12][1] ),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10214_ (.A1(_05053_),
    .A2(_05055_),
    .B(_05056_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10215_ (.I(_03712_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10216_ (.A1(_04220_),
    .A2(_05050_),
    .B1(_05048_),
    .B2(\stack[12][2] ),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10217_ (.A1(_05057_),
    .A2(_05055_),
    .B(_05058_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10218_ (.I(_03716_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10219_ (.A1(_04222_),
    .A2(_05050_),
    .B1(_05048_),
    .B2(\stack[12][3] ),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10220_ (.A1(_05059_),
    .A2(_05055_),
    .B(_05060_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10221_ (.I(_03721_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10222_ (.I(_05047_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10223_ (.A1(_04225_),
    .A2(_05045_),
    .B1(_05062_),
    .B2(\stack[12][4] ),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10224_ (.A1(_05061_),
    .A2(_05055_),
    .B(_05063_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10225_ (.I(_03728_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10226_ (.A1(_04227_),
    .A2(_05045_),
    .B1(_05062_),
    .B2(\stack[12][5] ),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10227_ (.A1(_05064_),
    .A2(_05054_),
    .B(_05065_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10228_ (.I(_01963_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_03847_),
    .A2(_04016_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10230_ (.I(_01124_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10231_ (.A1(_05068_),
    .A2(_05051_),
    .B1(_05062_),
    .B2(\stack[12][6] ),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10232_ (.A1(_05066_),
    .A2(_05067_),
    .B(_05069_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10233_ (.A1(_04206_),
    .A2(_05051_),
    .B1(_05062_),
    .B2(\stack[12][7] ),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10234_ (.A1(_04205_),
    .A2(_05067_),
    .B(_05070_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10235_ (.A1(_01640_),
    .A2(_03991_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10236_ (.I(_05071_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10237_ (.A1(_03635_),
    .A2(_03701_),
    .A3(_03994_),
    .A4(_03945_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10238_ (.I(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10239_ (.I(_01643_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10240_ (.A1(_01715_),
    .A2(_03990_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10241_ (.A1(_05075_),
    .A2(_05073_),
    .A3(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10242_ (.I(_05077_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10243_ (.A1(_01758_),
    .A2(_05074_),
    .B1(_05078_),
    .B2(\stack[14][0] ),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_03890_),
    .A2(_05072_),
    .B(_05079_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10245_ (.A1(_04218_),
    .A2(_05074_),
    .B1(_05078_),
    .B2(\stack[14][1] ),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10246_ (.A1(_05053_),
    .A2(_05072_),
    .B(_05080_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10247_ (.A1(_04220_),
    .A2(_05074_),
    .B1(_05078_),
    .B2(\stack[14][2] ),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10248_ (.A1(_05057_),
    .A2(_05072_),
    .B(_05081_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10249_ (.I(_05077_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10250_ (.A1(_04222_),
    .A2(_05074_),
    .B1(_05082_),
    .B2(\stack[14][3] ),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10251_ (.A1(_05059_),
    .A2(_05072_),
    .B(_05083_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10252_ (.A1(_04225_),
    .A2(_05073_),
    .B1(_05082_),
    .B2(\stack[14][4] ),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10253_ (.A1(_05061_),
    .A2(_05071_),
    .B(_05084_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10254_ (.A1(_04227_),
    .A2(_05073_),
    .B1(_05082_),
    .B2(\stack[14][5] ),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10255_ (.A1(_05064_),
    .A2(_05071_),
    .B(_05085_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10256_ (.A1(_01933_),
    .A2(_04016_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10257_ (.A1(\stack[14][6] ),
    .A2(_05078_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10258_ (.A1(_03908_),
    .A2(_05086_),
    .B1(_05071_),
    .B2(_03733_),
    .C(_05087_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10259_ (.A1(_04206_),
    .A2(_05076_),
    .B1(_05082_),
    .B2(\stack[14][7] ),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10260_ (.A1(_04205_),
    .A2(_05086_),
    .B(_05088_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10261_ (.A1(_01676_),
    .A2(_03701_),
    .A3(_03994_),
    .A4(_03945_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10262_ (.I(_05089_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10263_ (.A1(_03898_),
    .A2(_05090_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10264_ (.A1(_01638_),
    .A2(_03198_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10265_ (.I(_05092_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10266_ (.A1(_05075_),
    .A2(_05089_),
    .A3(_05092_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10267_ (.I(_05094_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10268_ (.A1(_04915_),
    .A2(_05093_),
    .B1(_05095_),
    .B2(\stack[30][0] ),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10269_ (.A1(_05091_),
    .A2(_05096_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10270_ (.I(_05093_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10271_ (.I(_05097_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10272_ (.A1(_01793_),
    .A2(_05090_),
    .B1(_05095_),
    .B2(\stack[30][1] ),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10273_ (.A1(_05053_),
    .A2(_05098_),
    .B(_05099_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10274_ (.A1(_01825_),
    .A2(_05090_),
    .B1(_05095_),
    .B2(\stack[30][2] ),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10275_ (.A1(_05057_),
    .A2(_05098_),
    .B(_05100_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10276_ (.I(_05094_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10277_ (.A1(_01857_),
    .A2(_05090_),
    .B1(_05101_),
    .B2(\stack[30][3] ),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10278_ (.A1(_05059_),
    .A2(_05098_),
    .B(_05102_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10279_ (.A1(_01888_),
    .A2(_05089_),
    .B1(_05101_),
    .B2(\stack[30][4] ),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10280_ (.A1(_05061_),
    .A2(_05098_),
    .B(_05103_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10281_ (.A1(_01923_),
    .A2(_05089_),
    .B1(_05101_),
    .B2(\stack[30][5] ),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10282_ (.A1(_05064_),
    .A2(_05097_),
    .B(_05104_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10283_ (.A1(_03909_),
    .A2(_03232_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10284_ (.A1(\stack[30][6] ),
    .A2(_05095_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10285_ (.A1(_03238_),
    .A2(_05093_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10286_ (.A1(_03908_),
    .A2(_05105_),
    .B(_05106_),
    .C(_05107_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10287_ (.A1(_04994_),
    .A2(_05093_),
    .B1(_05101_),
    .B2(\stack[30][7] ),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10288_ (.A1(_03854_),
    .A2(_05105_),
    .B(_05108_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10289_ (.A1(_03186_),
    .A2(_03188_),
    .A3(_03828_),
    .A4(_03702_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10290_ (.A1(_03743_),
    .A2(_03940_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10291_ (.A1(_03740_),
    .A2(_05109_),
    .A3(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10292_ (.I(_05111_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10293_ (.A1(\stack[27][0] ),
    .A2(_05112_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10294_ (.I(_05109_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10295_ (.I(_05110_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10296_ (.A1(_04191_),
    .A2(_05114_),
    .B1(_05115_),
    .B2(_04167_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10297_ (.A1(_05113_),
    .A2(_05116_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10298_ (.A1(_03870_),
    .A2(_03941_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10299_ (.I(_05111_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10300_ (.A1(\stack[27][1] ),
    .A2(_05118_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10301_ (.A1(_03752_),
    .A2(_05114_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10302_ (.A1(_03869_),
    .A2(_05117_),
    .B(_05119_),
    .C(_05120_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10303_ (.A1(\stack[27][2] ),
    .A2(_05112_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10304_ (.A1(_03218_),
    .A2(_05114_),
    .B1(_05115_),
    .B2(_04100_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10305_ (.A1(_05121_),
    .A2(_05122_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(\stack[27][3] ),
    .A2(_05112_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10307_ (.A1(_03221_),
    .A2(_05109_),
    .B1(_05115_),
    .B2(_04103_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10308_ (.A1(_05123_),
    .A2(_05124_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10309_ (.A1(\stack[27][4] ),
    .A2(_05118_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10310_ (.A1(_03762_),
    .A2(_05114_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10311_ (.A1(_03879_),
    .A2(_05117_),
    .B(_05125_),
    .C(_05126_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10312_ (.A1(_03228_),
    .A2(_05109_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10313_ (.A1(\stack[27][5] ),
    .A2(_05112_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10314_ (.A1(_03882_),
    .A2(_05117_),
    .B(_05127_),
    .C(_05128_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10315_ (.A1(_03663_),
    .A2(_03964_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10316_ (.A1(_05068_),
    .A2(_05115_),
    .B1(_05118_),
    .B2(\stack[27][6] ),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10317_ (.A1(_05066_),
    .A2(_05129_),
    .B(_05130_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(\stack[27][7] ),
    .A2(_05118_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10319_ (.A1(_04137_),
    .A2(_05129_),
    .B1(_05117_),
    .B2(_04112_),
    .C(_05131_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10320_ (.A1(_03858_),
    .A2(_04209_),
    .A3(_04026_),
    .A4(_03233_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10321_ (.A1(_03202_),
    .A2(_03643_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10322_ (.A1(_05075_),
    .A2(_05132_),
    .A3(_05133_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10323_ (.I(_05134_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10324_ (.A1(\stack[16][0] ),
    .A2(_05135_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10325_ (.I(_05132_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10326_ (.I(_05133_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10327_ (.A1(_04191_),
    .A2(_05137_),
    .B1(_05138_),
    .B2(_04915_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10328_ (.A1(_05136_),
    .A2(_05139_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10329_ (.I(_05138_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10330_ (.I(_05140_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10331_ (.A1(_01793_),
    .A2(_05137_),
    .B1(_05135_),
    .B2(\stack[16][1] ),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10332_ (.A1(_05053_),
    .A2(_05141_),
    .B(_05142_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10333_ (.A1(_01825_),
    .A2(_05137_),
    .B1(_05135_),
    .B2(\stack[16][2] ),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_05057_),
    .A2(_05141_),
    .B(_05143_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10335_ (.A1(_01857_),
    .A2(_05137_),
    .B1(_05135_),
    .B2(\stack[16][3] ),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10336_ (.A1(_05059_),
    .A2(_05141_),
    .B(_05144_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10337_ (.I(_05134_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10338_ (.A1(_01888_),
    .A2(_05132_),
    .B1(_05145_),
    .B2(\stack[16][4] ),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10339_ (.A1(_05061_),
    .A2(_05141_),
    .B(_05146_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10340_ (.A1(_01923_),
    .A2(_05132_),
    .B1(_05145_),
    .B2(\stack[16][5] ),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10341_ (.A1(_05064_),
    .A2(_05140_),
    .B(_05147_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10342_ (.A1(_03847_),
    .A2(_03662_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10343_ (.A1(_05068_),
    .A2(_05138_),
    .B1(_05145_),
    .B2(\stack[16][6] ),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10344_ (.A1(_05066_),
    .A2(_05148_),
    .B(_05149_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10345_ (.A1(_04994_),
    .A2(_05138_),
    .B1(_05145_),
    .B2(\stack[16][7] ),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10346_ (.A1(_03854_),
    .A2(_05148_),
    .B(_05150_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10347_ (.A1(_03668_),
    .A2(_01637_),
    .A3(_03630_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10348_ (.I(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10349_ (.A1(_03858_),
    .A2(_04209_),
    .A3(_03189_),
    .A4(_03690_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10350_ (.I(_05153_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10351_ (.A1(_03643_),
    .A2(_03996_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10352_ (.A1(_05075_),
    .A2(_05153_),
    .A3(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10353_ (.I(_05156_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10354_ (.A1(_01758_),
    .A2(_05154_),
    .B1(_05157_),
    .B2(\stack[17][0] ),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10355_ (.A1(_03890_),
    .A2(_05152_),
    .B(_05158_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10356_ (.A1(_01793_),
    .A2(_05154_),
    .B1(_05157_),
    .B2(\stack[17][1] ),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10357_ (.A1(_03869_),
    .A2(_05152_),
    .B(_05159_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10358_ (.A1(_01825_),
    .A2(_05154_),
    .B1(_05157_),
    .B2(\stack[17][2] ),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10359_ (.A1(_01796_),
    .A2(_05152_),
    .B(_05160_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10360_ (.I(_05156_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10361_ (.A1(_01857_),
    .A2(_05154_),
    .B1(_05161_),
    .B2(\stack[17][3] ),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10362_ (.A1(_01828_),
    .A2(_05152_),
    .B(_05162_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10363_ (.A1(_01888_),
    .A2(_05153_),
    .B1(_05161_),
    .B2(\stack[17][4] ),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10364_ (.A1(_03879_),
    .A2(_05151_),
    .B(_05163_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10365_ (.A1(_01923_),
    .A2(_05153_),
    .B1(_05161_),
    .B2(\stack[17][5] ),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10366_ (.A1(_03882_),
    .A2(_05151_),
    .B(_05164_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10367_ (.A1(_03662_),
    .A2(_03692_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10368_ (.A1(_05068_),
    .A2(_05155_),
    .B1(_05161_),
    .B2(\stack[17][6] ),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10369_ (.A1(_05066_),
    .A2(_05165_),
    .B(_05166_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10370_ (.A1(\stack[17][7] ),
    .A2(_05157_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10371_ (.A1(_04137_),
    .A2(_05165_),
    .B1(_05151_),
    .B2(_03855_),
    .C(_05167_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10372_ (.A1(_03858_),
    .A2(_03188_),
    .A3(_03189_),
    .A4(_03702_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10373_ (.A1(_03870_),
    .A2(_03991_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10374_ (.A1(_03261_),
    .A2(_05168_),
    .A3(_05169_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10375_ (.I(_05170_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10376_ (.I(_05168_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10377_ (.A1(_03633_),
    .A2(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10378_ (.I(_05169_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10379_ (.A1(_04915_),
    .A2(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10380_ (.A1(_01352_),
    .A2(_05171_),
    .B(_05173_),
    .C(_05175_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10381_ (.I(\stack[15][1] ),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10382_ (.A1(_03215_),
    .A2(_05172_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(net145),
    .A2(_05174_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10384_ (.A1(_05176_),
    .A2(_05171_),
    .B(_05177_),
    .C(_05178_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10385_ (.I(\stack[15][2] ),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10386_ (.A1(_03218_),
    .A2(_05172_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10387_ (.A1(_04100_),
    .A2(_05174_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10388_ (.A1(_05179_),
    .A2(_05171_),
    .B(_05180_),
    .C(_05181_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10389_ (.I(\stack[15][3] ),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10390_ (.I(_05168_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10391_ (.A1(_03221_),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10392_ (.A1(_04103_),
    .A2(_05174_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10393_ (.A1(_05182_),
    .A2(_05171_),
    .B(_05184_),
    .C(_05185_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10394_ (.I(\stack[15][4] ),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10395_ (.A1(_03224_),
    .A2(_05183_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10396_ (.I(_05169_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10397_ (.A1(net148),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10398_ (.A1(_05186_),
    .A2(_05170_),
    .B(_05187_),
    .C(_05189_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10399_ (.A1(_03724_),
    .A2(_05172_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10400_ (.A1(_04374_),
    .A2(_05183_),
    .A3(_05169_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10401_ (.A1(net149),
    .A2(_05188_),
    .B1(_05191_),
    .B2(\stack[15][5] ),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10402_ (.A1(_05190_),
    .A2(_05192_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10403_ (.I(_05183_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10404_ (.A1(_01125_),
    .A2(_05188_),
    .B1(_05191_),
    .B2(\stack[15][6] ),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10405_ (.A1(_03963_),
    .A2(_05193_),
    .B(_05194_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10406_ (.A1(_04994_),
    .A2(_05188_),
    .B1(_05191_),
    .B2(\stack[15][7] ),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10407_ (.A1(_03854_),
    .A2(_05193_),
    .B(_05195_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10408_ (.D(_00000_),
    .CLK(clknet_leaf_139_clock),
    .Q(\stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10409_ (.D(_00001_),
    .CLK(clknet_4_7_0_clock),
    .Q(\stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10410_ (.D(_00002_),
    .CLK(clknet_leaf_139_clock),
    .Q(\stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10411_ (.D(_00003_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10412_ (.D(_00004_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10413_ (.D(_00005_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10414_ (.D(_00006_),
    .CLK(clknet_4_3_0_clock),
    .Q(\stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10415_ (.D(_00007_),
    .CLK(clknet_leaf_3_clock),
    .Q(\stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10416_ (.D(_00008_),
    .CLK(clknet_leaf_40_clock),
    .Q(\mem.dff_data_ready ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10417_ (.D(_00009_),
    .CLK(clknet_leaf_39_clock),
    .Q(\mem.mem_dff.cycles[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10418_ (.D(_00010_),
    .CLK(clknet_leaf_39_clock),
    .Q(\mem.mem_dff.cycles[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10419_ (.D(_00011_),
    .CLK(clknet_leaf_122_clock),
    .Q(\mem.mem_dff.code_mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10420_ (.D(_00012_),
    .CLK(clknet_leaf_122_clock),
    .Q(\mem.mem_dff.code_mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10421_ (.D(_00013_),
    .CLK(clknet_leaf_122_clock),
    .Q(\mem.mem_dff.code_mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10422_ (.D(_00014_),
    .CLK(clknet_leaf_53_clock),
    .Q(\mem.mem_dff.code_mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10423_ (.D(_00015_),
    .CLK(clknet_leaf_54_clock),
    .Q(\mem.mem_dff.code_mem[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10424_ (.D(_00016_),
    .CLK(clknet_leaf_54_clock),
    .Q(\mem.mem_dff.code_mem[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10425_ (.D(_00017_),
    .CLK(clknet_leaf_54_clock),
    .Q(\mem.mem_dff.code_mem[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10426_ (.D(_00018_),
    .CLK(clknet_leaf_55_clock),
    .Q(\mem.mem_dff.code_mem[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10427_ (.D(_00019_),
    .CLK(clknet_leaf_60_clock),
    .Q(\mem.mem_dff.code_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10428_ (.D(_00020_),
    .CLK(clknet_leaf_61_clock),
    .Q(\mem.mem_dff.code_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10429_ (.D(_00021_),
    .CLK(clknet_leaf_61_clock),
    .Q(\mem.mem_dff.code_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10430_ (.D(_00022_),
    .CLK(clknet_leaf_75_clock),
    .Q(\mem.mem_dff.code_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10431_ (.D(_00023_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10432_ (.D(_00024_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10433_ (.D(_00025_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10434_ (.D(_00026_),
    .CLK(clknet_leaf_75_clock),
    .Q(\mem.mem_dff.code_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10435_ (.D(_00027_),
    .CLK(clknet_leaf_73_clock),
    .Q(\mem.mem_dff.code_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10436_ (.D(_00028_),
    .CLK(clknet_leaf_74_clock),
    .Q(\mem.mem_dff.code_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10437_ (.D(_00029_),
    .CLK(clknet_leaf_73_clock),
    .Q(\mem.mem_dff.code_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10438_ (.D(_00030_),
    .CLK(clknet_leaf_75_clock),
    .Q(\mem.mem_dff.code_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10439_ (.D(_00031_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10440_ (.D(_00032_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10441_ (.D(_00033_),
    .CLK(clknet_leaf_67_clock),
    .Q(\mem.mem_dff.code_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10442_ (.D(_00034_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10443_ (.D(_00035_),
    .CLK(clknet_leaf_74_clock),
    .Q(\mem.mem_dff.code_mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10444_ (.D(_00036_),
    .CLK(clknet_leaf_74_clock),
    .Q(\mem.mem_dff.code_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10445_ (.D(_00037_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10446_ (.D(_00038_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10447_ (.D(_00039_),
    .CLK(clknet_leaf_69_clock),
    .Q(\mem.mem_dff.code_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10448_ (.D(_00040_),
    .CLK(clknet_leaf_69_clock),
    .Q(\mem.mem_dff.code_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10449_ (.D(_00041_),
    .CLK(clknet_leaf_68_clock),
    .Q(\mem.mem_dff.code_mem[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10450_ (.D(_00042_),
    .CLK(clknet_leaf_69_clock),
    .Q(\mem.mem_dff.code_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10451_ (.D(_00043_),
    .CLK(clknet_leaf_73_clock),
    .Q(\mem.mem_dff.code_mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10452_ (.D(_00044_),
    .CLK(clknet_leaf_72_clock),
    .Q(\mem.mem_dff.code_mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10453_ (.D(_00045_),
    .CLK(clknet_leaf_73_clock),
    .Q(\mem.mem_dff.code_mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10454_ (.D(_00046_),
    .CLK(clknet_leaf_71_clock),
    .Q(\mem.mem_dff.code_mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10455_ (.D(_00047_),
    .CLK(clknet_leaf_70_clock),
    .Q(\mem.mem_dff.code_mem[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10456_ (.D(_00048_),
    .CLK(clknet_leaf_70_clock),
    .Q(\mem.mem_dff.code_mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10457_ (.D(_00049_),
    .CLK(clknet_leaf_70_clock),
    .Q(\mem.mem_dff.code_mem[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10458_ (.D(_00050_),
    .CLK(clknet_leaf_70_clock),
    .Q(\mem.mem_dff.code_mem[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10459_ (.D(_00051_),
    .CLK(clknet_leaf_72_clock),
    .Q(\mem.mem_dff.code_mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10460_ (.D(_00052_),
    .CLK(clknet_leaf_85_clock),
    .Q(\mem.mem_dff.code_mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10461_ (.D(_00053_),
    .CLK(clknet_leaf_72_clock),
    .Q(\mem.mem_dff.code_mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10462_ (.D(_00054_),
    .CLK(clknet_leaf_71_clock),
    .Q(\mem.mem_dff.code_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10463_ (.D(_00055_),
    .CLK(clknet_leaf_85_clock),
    .Q(\mem.mem_dff.code_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10464_ (.D(_00056_),
    .CLK(clknet_leaf_85_clock),
    .Q(\mem.mem_dff.code_mem[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10465_ (.D(_00057_),
    .CLK(clknet_leaf_70_clock),
    .Q(\mem.mem_dff.code_mem[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10466_ (.D(_00058_),
    .CLK(clknet_leaf_85_clock),
    .Q(\mem.mem_dff.code_mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10467_ (.D(_00059_),
    .CLK(clknet_leaf_57_clock),
    .Q(\mem.mem_dff.code_mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10468_ (.D(_00060_),
    .CLK(clknet_leaf_56_clock),
    .Q(\mem.mem_dff.code_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10469_ (.D(_00061_),
    .CLK(clknet_leaf_56_clock),
    .Q(\mem.mem_dff.code_mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10470_ (.D(_00062_),
    .CLK(clknet_leaf_57_clock),
    .Q(\mem.mem_dff.code_mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10471_ (.D(_00063_),
    .CLK(clknet_leaf_58_clock),
    .Q(\mem.mem_dff.code_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10472_ (.D(_00064_),
    .CLK(clknet_leaf_58_clock),
    .Q(\mem.mem_dff.code_mem[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10473_ (.D(_00065_),
    .CLK(clknet_leaf_58_clock),
    .Q(\mem.mem_dff.code_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10474_ (.D(_00066_),
    .CLK(clknet_leaf_57_clock),
    .Q(\mem.mem_dff.code_mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10475_ (.D(_00067_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10476_ (.D(_00068_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10477_ (.D(_00069_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10478_ (.D(_00070_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10479_ (.D(_00071_),
    .CLK(clknet_leaf_114_clock),
    .Q(\mem.mem_dff.code_mem[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10480_ (.D(_00072_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10481_ (.D(_00073_),
    .CLK(clknet_leaf_114_clock),
    .Q(\mem.mem_dff.code_mem[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10482_ (.D(_00074_),
    .CLK(clknet_leaf_123_clock),
    .Q(\mem.mem_dff.code_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10483_ (.D(_00075_),
    .CLK(clknet_leaf_56_clock),
    .Q(\mem.mem_dff.code_mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10484_ (.D(_00076_),
    .CLK(clknet_leaf_56_clock),
    .Q(\mem.mem_dff.code_mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10485_ (.D(_00077_),
    .CLK(clknet_leaf_56_clock),
    .Q(\mem.mem_dff.code_mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10486_ (.D(_00078_),
    .CLK(clknet_leaf_119_clock),
    .Q(\mem.mem_dff.code_mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10487_ (.D(_00079_),
    .CLK(clknet_leaf_118_clock),
    .Q(\mem.mem_dff.code_mem[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10488_ (.D(_00080_),
    .CLK(clknet_leaf_99_clock),
    .Q(\mem.mem_dff.code_mem[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10489_ (.D(_00081_),
    .CLK(clknet_leaf_118_clock),
    .Q(\mem.mem_dff.code_mem[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10490_ (.D(_00082_),
    .CLK(clknet_leaf_118_clock),
    .Q(\mem.mem_dff.code_mem[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10491_ (.D(_00083_),
    .CLK(clknet_leaf_120_clock),
    .Q(\mem.mem_dff.code_mem[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10492_ (.D(_00084_),
    .CLK(clknet_leaf_120_clock),
    .Q(\mem.mem_dff.code_mem[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10493_ (.D(_00085_),
    .CLK(clknet_leaf_120_clock),
    .Q(\mem.mem_dff.code_mem[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10494_ (.D(_00086_),
    .CLK(clknet_leaf_120_clock),
    .Q(\mem.mem_dff.code_mem[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10495_ (.D(_00087_),
    .CLK(clknet_leaf_117_clock),
    .Q(\mem.mem_dff.code_mem[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10496_ (.D(_00088_),
    .CLK(clknet_leaf_116_clock),
    .Q(\mem.mem_dff.code_mem[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10497_ (.D(_00089_),
    .CLK(clknet_leaf_117_clock),
    .Q(\mem.mem_dff.code_mem[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10498_ (.D(_00090_),
    .CLK(clknet_leaf_117_clock),
    .Q(\mem.mem_dff.code_mem[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10499_ (.D(_00091_),
    .CLK(clknet_leaf_108_clock),
    .Q(\mem.mem_dff.code_mem[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10500_ (.D(_00092_),
    .CLK(clknet_leaf_108_clock),
    .Q(\mem.mem_dff.code_mem[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10501_ (.D(_00093_),
    .CLK(clknet_leaf_108_clock),
    .Q(\mem.mem_dff.code_mem[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10502_ (.D(_00094_),
    .CLK(clknet_leaf_108_clock),
    .Q(\mem.mem_dff.code_mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10503_ (.D(_00095_),
    .CLK(clknet_leaf_107_clock),
    .Q(\mem.mem_dff.code_mem[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10504_ (.D(_00096_),
    .CLK(clknet_leaf_109_clock),
    .Q(\mem.mem_dff.code_mem[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10505_ (.D(_00097_),
    .CLK(clknet_leaf_106_clock),
    .Q(\mem.mem_dff.code_mem[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10506_ (.D(_00098_),
    .CLK(clknet_leaf_109_clock),
    .Q(\mem.mem_dff.code_mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10507_ (.D(_00099_),
    .CLK(clknet_leaf_111_clock),
    .Q(\mem.mem_dff.code_mem[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10508_ (.D(_00100_),
    .CLK(clknet_leaf_108_clock),
    .Q(\mem.mem_dff.code_mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10509_ (.D(_00101_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10510_ (.D(_00102_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10511_ (.D(_00103_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10512_ (.D(_00104_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10513_ (.D(_00105_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10514_ (.D(_00106_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10515_ (.D(_00107_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10516_ (.D(_00108_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10517_ (.D(_00109_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10518_ (.D(_00110_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10519_ (.D(_00111_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10520_ (.D(_00112_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10521_ (.D(_00113_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10522_ (.D(_00114_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10523_ (.D(_00115_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10524_ (.D(_00116_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10525_ (.D(_00117_),
    .CLK(clknet_leaf_110_clock),
    .Q(\mem.mem_dff.code_mem[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10526_ (.D(_00118_),
    .CLK(clknet_leaf_111_clock),
    .Q(\mem.mem_dff.code_mem[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10527_ (.D(_00119_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10528_ (.D(_00120_),
    .CLK(clknet_leaf_113_clock),
    .Q(\mem.mem_dff.code_mem[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10529_ (.D(_00121_),
    .CLK(clknet_leaf_113_clock),
    .Q(\mem.mem_dff.code_mem[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10530_ (.D(_00122_),
    .CLK(clknet_leaf_112_clock),
    .Q(\mem.mem_dff.code_mem[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10531_ (.D(_00123_),
    .CLK(clknet_leaf_124_clock),
    .Q(\mem.mem_dff.code_mem[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10532_ (.D(_00124_),
    .CLK(clknet_leaf_124_clock),
    .Q(\mem.mem_dff.code_mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10533_ (.D(_00125_),
    .CLK(clknet_leaf_124_clock),
    .Q(\mem.mem_dff.code_mem[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10534_ (.D(_00126_),
    .CLK(clknet_leaf_113_clock),
    .Q(\mem.mem_dff.code_mem[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10535_ (.D(_00127_),
    .CLK(clknet_leaf_114_clock),
    .Q(\mem.mem_dff.code_mem[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10536_ (.D(_00128_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10537_ (.D(_00129_),
    .CLK(clknet_leaf_113_clock),
    .Q(\mem.mem_dff.code_mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10538_ (.D(_00130_),
    .CLK(clknet_leaf_113_clock),
    .Q(\mem.mem_dff.code_mem[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10539_ (.D(_00131_),
    .CLK(clknet_leaf_98_clock),
    .Q(\mem.mem_dff.code_mem[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10540_ (.D(_00132_),
    .CLK(clknet_leaf_98_clock),
    .Q(\mem.mem_dff.code_mem[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10541_ (.D(_00133_),
    .CLK(clknet_leaf_97_clock),
    .Q(\mem.mem_dff.code_mem[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10542_ (.D(_00134_),
    .CLK(clknet_leaf_97_clock),
    .Q(\mem.mem_dff.code_mem[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10543_ (.D(_00135_),
    .CLK(clknet_leaf_97_clock),
    .Q(\mem.mem_dff.code_mem[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10544_ (.D(_00136_),
    .CLK(clknet_leaf_97_clock),
    .Q(\mem.mem_dff.code_mem[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10545_ (.D(_00137_),
    .CLK(clknet_leaf_96_clock),
    .Q(\mem.mem_dff.code_mem[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10546_ (.D(_00138_),
    .CLK(clknet_leaf_79_clock),
    .Q(\mem.mem_dff.code_mem[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10547_ (.D(_00139_),
    .CLK(clknet_leaf_79_clock),
    .Q(\mem.mem_dff.code_mem[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10548_ (.D(_00140_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10549_ (.D(_00141_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10550_ (.D(_00142_),
    .CLK(clknet_leaf_76_clock),
    .Q(\mem.mem_dff.code_mem[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10551_ (.D(_00143_),
    .CLK(clknet_leaf_79_clock),
    .Q(\mem.mem_dff.code_mem[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10552_ (.D(_00144_),
    .CLK(clknet_leaf_79_clock),
    .Q(\mem.mem_dff.code_mem[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10553_ (.D(_00145_),
    .CLK(clknet_leaf_80_clock),
    .Q(\mem.mem_dff.code_mem[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10554_ (.D(_00146_),
    .CLK(clknet_leaf_80_clock),
    .Q(\mem.mem_dff.code_mem[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10555_ (.D(_00147_),
    .CLK(clknet_leaf_95_clock),
    .Q(\mem.mem_dff.code_mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10556_ (.D(_00148_),
    .CLK(clknet_leaf_91_clock),
    .Q(\mem.mem_dff.code_mem[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10557_ (.D(_00149_),
    .CLK(clknet_leaf_91_clock),
    .Q(\mem.mem_dff.code_mem[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10558_ (.D(_00150_),
    .CLK(clknet_leaf_91_clock),
    .Q(\mem.mem_dff.code_mem[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10559_ (.D(_00151_),
    .CLK(clknet_leaf_96_clock),
    .Q(\mem.mem_dff.code_mem[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10560_ (.D(_00152_),
    .CLK(clknet_leaf_96_clock),
    .Q(\mem.mem_dff.code_mem[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10561_ (.D(_00153_),
    .CLK(clknet_leaf_96_clock),
    .Q(\mem.mem_dff.code_mem[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10562_ (.D(_00154_),
    .CLK(clknet_leaf_80_clock),
    .Q(\mem.mem_dff.code_mem[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10563_ (.D(_00155_),
    .CLK(clknet_4_15_0_clock),
    .Q(\mem.mem_dff.code_mem[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10564_ (.D(_00156_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10565_ (.D(_00157_),
    .CLK(clknet_leaf_73_clock),
    .Q(\mem.mem_dff.code_mem[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10566_ (.D(_00158_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10567_ (.D(_00159_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10568_ (.D(_00160_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10569_ (.D(_00161_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10570_ (.D(_00162_),
    .CLK(clknet_leaf_82_clock),
    .Q(\mem.mem_dff.code_mem[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10571_ (.D(_00163_),
    .CLK(clknet_leaf_81_clock),
    .Q(\mem.mem_dff.code_mem[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10572_ (.D(_00164_),
    .CLK(clknet_leaf_81_clock),
    .Q(\mem.mem_dff.code_mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10573_ (.D(_00165_),
    .CLK(clknet_leaf_81_clock),
    .Q(\mem.mem_dff.code_mem[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10574_ (.D(_00166_),
    .CLK(clknet_leaf_89_clock),
    .Q(\mem.mem_dff.code_mem[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10575_ (.D(_00167_),
    .CLK(clknet_leaf_89_clock),
    .Q(\mem.mem_dff.code_mem[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10576_ (.D(_00168_),
    .CLK(clknet_leaf_90_clock),
    .Q(\mem.mem_dff.code_mem[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10577_ (.D(_00169_),
    .CLK(clknet_leaf_91_clock),
    .Q(\mem.mem_dff.code_mem[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10578_ (.D(_00170_),
    .CLK(clknet_leaf_89_clock),
    .Q(\mem.mem_dff.code_mem[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10579_ (.D(_00171_),
    .CLK(clknet_leaf_84_clock),
    .Q(\mem.mem_dff.code_mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10580_ (.D(_00172_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10581_ (.D(_00173_),
    .CLK(clknet_leaf_84_clock),
    .Q(\mem.mem_dff.code_mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10582_ (.D(_00174_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10583_ (.D(_00175_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10584_ (.D(_00176_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10585_ (.D(_00177_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10586_ (.D(_00178_),
    .CLK(clknet_leaf_86_clock),
    .Q(\mem.mem_dff.code_mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10587_ (.D(_00179_),
    .CLK(clknet_leaf_81_clock),
    .Q(\mem.mem_dff.code_mem[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10588_ (.D(_00180_),
    .CLK(clknet_leaf_88_clock),
    .Q(\mem.mem_dff.code_mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10589_ (.D(_00181_),
    .CLK(clknet_leaf_88_clock),
    .Q(\mem.mem_dff.code_mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10590_ (.D(_00182_),
    .CLK(clknet_leaf_87_clock),
    .Q(\mem.mem_dff.code_mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10591_ (.D(_00183_),
    .CLK(clknet_leaf_87_clock),
    .Q(\mem.mem_dff.code_mem[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10592_ (.D(_00184_),
    .CLK(clknet_leaf_87_clock),
    .Q(\mem.mem_dff.code_mem[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10593_ (.D(_00185_),
    .CLK(clknet_leaf_87_clock),
    .Q(\mem.mem_dff.code_mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10594_ (.D(_00186_),
    .CLK(clknet_leaf_90_clock),
    .Q(\mem.mem_dff.code_mem[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10595_ (.D(_00187_),
    .CLK(clknet_leaf_99_clock),
    .Q(\mem.mem_dff.code_mem[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10596_ (.D(_00188_),
    .CLK(clknet_leaf_99_clock),
    .Q(\mem.mem_dff.code_mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10597_ (.D(_00189_),
    .CLK(clknet_leaf_99_clock),
    .Q(\mem.mem_dff.code_mem[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10598_ (.D(_00190_),
    .CLK(clknet_leaf_99_clock),
    .Q(\mem.mem_dff.code_mem[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10599_ (.D(_00191_),
    .CLK(clknet_leaf_100_clock),
    .Q(\mem.mem_dff.code_mem[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10600_ (.D(_00192_),
    .CLK(clknet_leaf_100_clock),
    .Q(\mem.mem_dff.code_mem[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10601_ (.D(_00193_),
    .CLK(clknet_leaf_100_clock),
    .Q(\mem.mem_dff.code_mem[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10602_ (.D(_00194_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10603_ (.D(_00195_),
    .CLK(clknet_leaf_93_clock),
    .Q(\mem.mem_dff.code_mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10604_ (.D(_00196_),
    .CLK(clknet_leaf_93_clock),
    .Q(\mem.mem_dff.code_mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10605_ (.D(_00197_),
    .CLK(clknet_leaf_93_clock),
    .Q(\mem.mem_dff.code_mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10606_ (.D(_00198_),
    .CLK(clknet_leaf_92_clock),
    .Q(\mem.mem_dff.code_mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10607_ (.D(_00199_),
    .CLK(clknet_leaf_92_clock),
    .Q(\mem.mem_dff.code_mem[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10608_ (.D(_00200_),
    .CLK(clknet_leaf_92_clock),
    .Q(\mem.mem_dff.code_mem[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10609_ (.D(_00201_),
    .CLK(clknet_leaf_92_clock),
    .Q(\mem.mem_dff.code_mem[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10610_ (.D(_00202_),
    .CLK(clknet_leaf_92_clock),
    .Q(\mem.mem_dff.code_mem[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10611_ (.D(_00203_),
    .CLK(clknet_leaf_107_clock),
    .Q(\mem.mem_dff.code_mem[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10612_ (.D(_00204_),
    .CLK(clknet_leaf_106_clock),
    .Q(\mem.mem_dff.code_mem[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10613_ (.D(_00205_),
    .CLK(clknet_leaf_106_clock),
    .Q(\mem.mem_dff.code_mem[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10614_ (.D(_00206_),
    .CLK(clknet_leaf_107_clock),
    .Q(\mem.mem_dff.code_mem[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10615_ (.D(_00207_),
    .CLK(clknet_leaf_106_clock),
    .Q(\mem.mem_dff.code_mem[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10616_ (.D(_00208_),
    .CLK(clknet_leaf_105_clock),
    .Q(\mem.mem_dff.code_mem[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10617_ (.D(_00209_),
    .CLK(clknet_leaf_106_clock),
    .Q(\mem.mem_dff.code_mem[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10618_ (.D(_00210_),
    .CLK(clknet_leaf_105_clock),
    .Q(\mem.mem_dff.code_mem[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10619_ (.D(_00211_),
    .CLK(clknet_leaf_105_clock),
    .Q(\mem.mem_dff.code_mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10620_ (.D(_00212_),
    .CLK(clknet_leaf_105_clock),
    .Q(\mem.mem_dff.code_mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10621_ (.D(_00213_),
    .CLK(clknet_leaf_105_clock),
    .Q(\mem.mem_dff.code_mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10622_ (.D(_00214_),
    .CLK(clknet_leaf_104_clock),
    .Q(\mem.mem_dff.code_mem[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10623_ (.D(_00215_),
    .CLK(clknet_leaf_104_clock),
    .Q(\mem.mem_dff.code_mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10624_ (.D(_00216_),
    .CLK(clknet_leaf_104_clock),
    .Q(\mem.mem_dff.code_mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10625_ (.D(_00217_),
    .CLK(clknet_leaf_104_clock),
    .Q(\mem.mem_dff.code_mem[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10626_ (.D(_00218_),
    .CLK(clknet_leaf_104_clock),
    .Q(\mem.mem_dff.code_mem[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10627_ (.D(_00219_),
    .CLK(clknet_leaf_101_clock),
    .Q(\mem.mem_dff.code_mem[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10628_ (.D(_00220_),
    .CLK(clknet_leaf_102_clock),
    .Q(\mem.mem_dff.code_mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10629_ (.D(_00221_),
    .CLK(clknet_leaf_102_clock),
    .Q(\mem.mem_dff.code_mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10630_ (.D(_00222_),
    .CLK(clknet_leaf_102_clock),
    .Q(\mem.mem_dff.code_mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10631_ (.D(_00223_),
    .CLK(clknet_leaf_101_clock),
    .Q(\mem.mem_dff.code_mem[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10632_ (.D(_00224_),
    .CLK(clknet_leaf_115_clock),
    .Q(\mem.mem_dff.code_mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10633_ (.D(_00225_),
    .CLK(clknet_leaf_101_clock),
    .Q(\mem.mem_dff.code_mem[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10634_ (.D(_00226_),
    .CLK(clknet_leaf_101_clock),
    .Q(\mem.mem_dff.code_mem[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10635_ (.D(_00227_),
    .CLK(clknet_leaf_100_clock),
    .Q(\mem.mem_dff.code_mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10636_ (.D(_00228_),
    .CLK(clknet_leaf_102_clock),
    .Q(\mem.mem_dff.code_mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10637_ (.D(_00229_),
    .CLK(clknet_leaf_102_clock),
    .Q(\mem.mem_dff.code_mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10638_ (.D(_00230_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10639_ (.D(_00231_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10640_ (.D(_00232_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10641_ (.D(_00233_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10642_ (.D(_00234_),
    .CLK(clknet_leaf_103_clock),
    .Q(\mem.mem_dff.code_mem[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10643_ (.D(_00235_),
    .CLK(clknet_leaf_120_clock),
    .Q(\mem.mem_dff.code_mem[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10644_ (.D(_00236_),
    .CLK(clknet_leaf_119_clock),
    .Q(\mem.mem_dff.code_mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10645_ (.D(_00237_),
    .CLK(clknet_4_12_0_clock),
    .Q(\mem.mem_dff.code_mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10646_ (.D(_00238_),
    .CLK(clknet_leaf_117_clock),
    .Q(\mem.mem_dff.code_mem[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10647_ (.D(_00239_),
    .CLK(clknet_leaf_116_clock),
    .Q(\mem.mem_dff.code_mem[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10648_ (.D(_00240_),
    .CLK(clknet_leaf_116_clock),
    .Q(\mem.mem_dff.code_mem[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10649_ (.D(_00241_),
    .CLK(clknet_leaf_116_clock),
    .Q(\mem.mem_dff.code_mem[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10650_ (.D(_00242_),
    .CLK(clknet_leaf_101_clock),
    .Q(\mem.mem_dff.code_mem[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10651_ (.D(_00243_),
    .CLK(clknet_leaf_94_clock),
    .Q(\mem.mem_dff.code_mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10652_ (.D(_00244_),
    .CLK(clknet_leaf_94_clock),
    .Q(\mem.mem_dff.code_mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10653_ (.D(_00245_),
    .CLK(clknet_leaf_94_clock),
    .Q(\mem.mem_dff.code_mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10654_ (.D(_00246_),
    .CLK(clknet_leaf_94_clock),
    .Q(\mem.mem_dff.code_mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10655_ (.D(_00247_),
    .CLK(clknet_leaf_95_clock),
    .Q(\mem.mem_dff.code_mem[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10656_ (.D(_00248_),
    .CLK(clknet_leaf_95_clock),
    .Q(\mem.mem_dff.code_mem[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10657_ (.D(_00249_),
    .CLK(clknet_leaf_95_clock),
    .Q(\mem.mem_dff.code_mem[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10658_ (.D(_00250_),
    .CLK(clknet_leaf_93_clock),
    .Q(\mem.mem_dff.code_mem[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10659_ (.D(_00251_),
    .CLK(clknet_leaf_78_clock),
    .Q(\mem.mem_dff.code_mem[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10660_ (.D(_00252_),
    .CLK(clknet_leaf_78_clock),
    .Q(\mem.mem_dff.code_mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10661_ (.D(_00253_),
    .CLK(clknet_leaf_57_clock),
    .Q(\mem.mem_dff.code_mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10662_ (.D(_00254_),
    .CLK(clknet_leaf_78_clock),
    .Q(\mem.mem_dff.code_mem[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10663_ (.D(_00255_),
    .CLK(clknet_leaf_77_clock),
    .Q(\mem.mem_dff.code_mem[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10664_ (.D(_00256_),
    .CLK(clknet_leaf_77_clock),
    .Q(\mem.mem_dff.code_mem[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10665_ (.D(_00257_),
    .CLK(clknet_leaf_77_clock),
    .Q(\mem.mem_dff.code_mem[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10666_ (.D(_00258_),
    .CLK(clknet_leaf_57_clock),
    .Q(\mem.mem_dff.code_mem[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10667_ (.D(_00259_),
    .CLK(clknet_leaf_55_clock),
    .Q(\mem.mem_dff.code_mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10668_ (.D(_00260_),
    .CLK(clknet_leaf_55_clock),
    .Q(\mem.mem_dff.code_mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10669_ (.D(_00261_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.code_mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10670_ (.D(_00262_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.code_mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10671_ (.D(_00263_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.code_mem[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10672_ (.D(_00264_),
    .CLK(clknet_leaf_60_clock),
    .Q(\mem.mem_dff.code_mem[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10673_ (.D(_00265_),
    .CLK(clknet_leaf_60_clock),
    .Q(\mem.mem_dff.code_mem[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10674_ (.D(_00266_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.code_mem[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10675_ (.D(_00267_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.mem_dff.data_mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10676_ (.D(_00268_),
    .CLK(clknet_leaf_48_clock),
    .Q(\mem.mem_dff.data_mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10677_ (.D(_00269_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.mem_dff.data_mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10678_ (.D(_00270_),
    .CLK(clknet_4_9_0_clock),
    .Q(\mem.mem_dff.data_mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10679_ (.D(_00271_),
    .CLK(clknet_leaf_51_clock),
    .Q(\mem.mem_dff.data_mem[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10680_ (.D(_00272_),
    .CLK(clknet_leaf_51_clock),
    .Q(\mem.mem_dff.data_mem[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10681_ (.D(_00273_),
    .CLK(clknet_leaf_51_clock),
    .Q(\mem.mem_dff.data_mem[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10682_ (.D(_00274_),
    .CLK(clknet_leaf_54_clock),
    .Q(\mem.mem_dff.data_mem[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10683_ (.D(_00275_),
    .CLK(clknet_leaf_60_clock),
    .Q(\mem.mem_dff.data_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10684_ (.D(_00276_),
    .CLK(clknet_leaf_62_clock),
    .Q(\mem.mem_dff.data_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10685_ (.D(_00277_),
    .CLK(clknet_leaf_60_clock),
    .Q(\mem.mem_dff.data_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10686_ (.D(_00278_),
    .CLK(clknet_leaf_62_clock),
    .Q(\mem.mem_dff.data_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10687_ (.D(_00279_),
    .CLK(clknet_leaf_61_clock),
    .Q(\mem.mem_dff.data_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10688_ (.D(_00280_),
    .CLK(clknet_leaf_61_clock),
    .Q(\mem.mem_dff.data_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10689_ (.D(_00281_),
    .CLK(clknet_leaf_67_clock),
    .Q(\mem.mem_dff.data_mem[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10690_ (.D(_00282_),
    .CLK(clknet_leaf_61_clock),
    .Q(\mem.mem_dff.data_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10691_ (.D(_00283_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.data_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10692_ (.D(_00284_),
    .CLK(clknet_leaf_55_clock),
    .Q(\mem.mem_dff.data_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10693_ (.D(_00285_),
    .CLK(clknet_leaf_54_clock),
    .Q(\mem.mem_dff.data_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10694_ (.D(_00286_),
    .CLK(clknet_4_14_0_clock),
    .Q(\mem.mem_dff.data_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10695_ (.D(_00287_),
    .CLK(clknet_leaf_62_clock),
    .Q(\mem.mem_dff.data_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10696_ (.D(_00288_),
    .CLK(clknet_leaf_59_clock),
    .Q(\mem.mem_dff.data_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10697_ (.D(_00289_),
    .CLK(clknet_leaf_62_clock),
    .Q(\mem.mem_dff.data_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10698_ (.D(_00290_),
    .CLK(clknet_leaf_62_clock),
    .Q(\mem.mem_dff.data_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10699_ (.D(_00291_),
    .CLK(clknet_leaf_66_clock),
    .Q(\mem.mem_dff.data_mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10700_ (.D(_00292_),
    .CLK(clknet_leaf_66_clock),
    .Q(\mem.mem_dff.data_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10701_ (.D(_00293_),
    .CLK(clknet_leaf_66_clock),
    .Q(\mem.mem_dff.data_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10702_ (.D(_00294_),
    .CLK(clknet_leaf_66_clock),
    .Q(\mem.mem_dff.data_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10703_ (.D(_00295_),
    .CLK(clknet_leaf_66_clock),
    .Q(\mem.mem_dff.data_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10704_ (.D(_00296_),
    .CLK(clknet_leaf_29_clock),
    .Q(\mem.mem_dff.data_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10705_ (.D(_00297_),
    .CLK(clknet_leaf_65_clock),
    .Q(\mem.mem_dff.data_mem[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10706_ (.D(_00298_),
    .CLK(clknet_leaf_29_clock),
    .Q(\mem.mem_dff.data_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10707_ (.D(_00299_),
    .CLK(clknet_leaf_30_clock),
    .Q(\mem.mem_dff.data_mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10708_ (.D(_00300_),
    .CLK(clknet_leaf_37_clock),
    .Q(\mem.mem_dff.data_mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10709_ (.D(_00301_),
    .CLK(clknet_leaf_37_clock),
    .Q(\mem.mem_dff.data_mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10710_ (.D(_00302_),
    .CLK(clknet_leaf_36_clock),
    .Q(\mem.mem_dff.data_mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10711_ (.D(_00303_),
    .CLK(clknet_leaf_30_clock),
    .Q(\mem.mem_dff.data_mem[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10712_ (.D(_00304_),
    .CLK(clknet_leaf_29_clock),
    .Q(\mem.mem_dff.data_mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10713_ (.D(_00305_),
    .CLK(clknet_leaf_29_clock),
    .Q(\mem.mem_dff.data_mem[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10714_ (.D(_00306_),
    .CLK(clknet_leaf_30_clock),
    .Q(\mem.mem_dff.data_mem[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10715_ (.D(_00307_),
    .CLK(clknet_leaf_31_clock),
    .Q(\mem.mem_dff.data_mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10716_ (.D(_00308_),
    .CLK(clknet_leaf_36_clock),
    .Q(\mem.mem_dff.data_mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10717_ (.D(_00309_),
    .CLK(clknet_leaf_36_clock),
    .Q(\mem.mem_dff.data_mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10718_ (.D(_00310_),
    .CLK(clknet_leaf_36_clock),
    .Q(\mem.mem_dff.data_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10719_ (.D(_00311_),
    .CLK(clknet_leaf_30_clock),
    .Q(\mem.mem_dff.data_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10720_ (.D(_00312_),
    .CLK(clknet_leaf_31_clock),
    .Q(\mem.mem_dff.data_mem[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10721_ (.D(_00313_),
    .CLK(clknet_leaf_29_clock),
    .Q(\mem.mem_dff.data_mem[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10722_ (.D(_00314_),
    .CLK(clknet_leaf_30_clock),
    .Q(\mem.mem_dff.data_mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10723_ (.D(_00315_),
    .CLK(clknet_leaf_50_clock),
    .Q(\mem.mem_dff.data_mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10724_ (.D(_00316_),
    .CLK(clknet_leaf_51_clock),
    .Q(\mem.mem_dff.data_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10725_ (.D(_00317_),
    .CLK(clknet_leaf_50_clock),
    .Q(\mem.mem_dff.data_mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10726_ (.D(_00318_),
    .CLK(clknet_leaf_51_clock),
    .Q(\mem.mem_dff.data_mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10727_ (.D(_00319_),
    .CLK(clknet_leaf_64_clock),
    .Q(\mem.mem_dff.data_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10728_ (.D(_00320_),
    .CLK(clknet_leaf_64_clock),
    .Q(\mem.mem_dff.data_mem[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10729_ (.D(_00321_),
    .CLK(clknet_leaf_64_clock),
    .Q(\mem.mem_dff.data_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10730_ (.D(_00322_),
    .CLK(clknet_leaf_64_clock),
    .Q(\mem.mem_dff.data_mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10731_ (.D(_00323_),
    .CLK(clknet_leaf_50_clock),
    .Q(\mem.mem_dff.data_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10732_ (.D(_00324_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.mem_dff.data_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10733_ (.D(_00325_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.mem_dff.data_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10734_ (.D(_00326_),
    .CLK(clknet_leaf_50_clock),
    .Q(\mem.mem_dff.data_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10735_ (.D(_00327_),
    .CLK(clknet_leaf_64_clock),
    .Q(\mem.mem_dff.data_mem[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10736_ (.D(_00328_),
    .CLK(clknet_leaf_65_clock),
    .Q(\mem.mem_dff.data_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10737_ (.D(_00329_),
    .CLK(clknet_leaf_65_clock),
    .Q(\mem.mem_dff.data_mem[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10738_ (.D(_00330_),
    .CLK(clknet_leaf_65_clock),
    .Q(\mem.mem_dff.data_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10739_ (.D(_00331_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10740_ (.D(_00332_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10741_ (.D(_00333_),
    .CLK(clknet_leaf_134_clock),
    .Q(\stack[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10742_ (.D(_00334_),
    .CLK(clknet_leaf_163_clock),
    .Q(\stack[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10743_ (.D(_00335_),
    .CLK(clknet_leaf_167_clock),
    .Q(\stack[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10744_ (.D(_00336_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10745_ (.D(_00337_),
    .CLK(clknet_leaf_3_clock),
    .Q(\stack[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10746_ (.D(_00338_),
    .CLK(clknet_leaf_3_clock),
    .Q(\stack[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10747_ (.D(_00339_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10748_ (.D(_00340_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10749_ (.D(_00341_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10750_ (.D(_00342_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10751_ (.D(_00343_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10752_ (.D(_00344_),
    .CLK(clknet_leaf_38_clock),
    .Q(\mem.io_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10753_ (.D(_00345_),
    .CLK(clknet_leaf_41_clock),
    .Q(\mem.io_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10754_ (.D(_00346_),
    .CLK(clknet_leaf_42_clock),
    .Q(\mem.io_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10755_ (.D(_00347_),
    .CLK(clknet_leaf_48_clock),
    .Q(\mem.dff_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10756_ (.D(_00348_),
    .CLK(clknet_leaf_48_clock),
    .Q(\mem.dff_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10757_ (.D(_00349_),
    .CLK(clknet_leaf_47_clock),
    .Q(\mem.dff_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10758_ (.D(_00350_),
    .CLK(clknet_leaf_47_clock),
    .Q(\mem.dff_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10759_ (.D(_00351_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.dff_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10760_ (.D(_00352_),
    .CLK(clknet_leaf_48_clock),
    .Q(\mem.dff_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10761_ (.D(_00353_),
    .CLK(clknet_leaf_37_clock),
    .Q(\mem.dff_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10762_ (.D(_00354_),
    .CLK(clknet_leaf_49_clock),
    .Q(\mem.dff_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10763_ (.D(_00355_),
    .CLK(clknet_leaf_37_clock),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10764_ (.D(_00356_),
    .CLK(clknet_leaf_37_clock),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10765_ (.D(_00357_),
    .CLK(clknet_leaf_37_clock),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10766_ (.D(_00358_),
    .CLK(clknet_leaf_36_clock),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10767_ (.D(_00359_),
    .CLK(clknet_leaf_31_clock),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10768_ (.D(_00360_),
    .CLK(clknet_leaf_31_clock),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10769_ (.D(_00361_),
    .CLK(clknet_leaf_31_clock),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10770_ (.D(_00362_),
    .CLK(clknet_leaf_31_clock),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10771_ (.D(_00363_),
    .CLK(clknet_leaf_53_clock),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10772_ (.D(_00364_),
    .CLK(clknet_leaf_53_clock),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10773_ (.D(_00365_),
    .CLK(clknet_leaf_53_clock),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10774_ (.D(_00366_),
    .CLK(clknet_leaf_53_clock),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10775_ (.D(_00367_),
    .CLK(clknet_leaf_122_clock),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10776_ (.D(_00368_),
    .CLK(clknet_leaf_122_clock),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10777_ (.D(_00369_),
    .CLK(clknet_leaf_53_clock),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10778_ (.D(_00370_),
    .CLK(clknet_leaf_122_clock),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10779_ (.D(_00371_),
    .CLK(clknet_leaf_41_clock),
    .Q(\mem.io_data_ready ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10780_ (.D(_00372_),
    .CLK(clknet_leaf_10_clock),
    .Q(\intr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10781_ (.D(_00373_),
    .CLK(clknet_leaf_135_clock),
    .Q(\stack[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10782_ (.D(_00374_),
    .CLK(clknet_leaf_135_clock),
    .Q(\stack[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10783_ (.D(_00375_),
    .CLK(clknet_leaf_135_clock),
    .Q(\stack[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10784_ (.D(_00376_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10785_ (.D(_00377_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10786_ (.D(_00378_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10787_ (.D(_00379_),
    .CLK(clknet_leaf_3_clock),
    .Q(\stack[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10788_ (.D(_00380_),
    .CLK(clknet_leaf_3_clock),
    .Q(\stack[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10789_ (.D(_00381_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10790_ (.D(_00382_),
    .CLK(clknet_leaf_135_clock),
    .Q(\stack[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10791_ (.D(_00383_),
    .CLK(clknet_leaf_135_clock),
    .Q(\stack[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10792_ (.D(_00384_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10793_ (.D(_00385_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10794_ (.D(_00386_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10795_ (.D(_00387_),
    .CLK(clknet_leaf_5_clock),
    .Q(\stack[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10796_ (.D(_00388_),
    .CLK(clknet_4_0_0_clock),
    .Q(\stack[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10797_ (.D(_00389_),
    .CLK(clknet_leaf_134_clock),
    .Q(\stack[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10798_ (.D(_00390_),
    .CLK(clknet_leaf_163_clock),
    .Q(\stack[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10799_ (.D(_00391_),
    .CLK(clknet_leaf_134_clock),
    .Q(\stack[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10800_ (.D(_00392_),
    .CLK(clknet_leaf_163_clock),
    .Q(\stack[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10801_ (.D(_00393_),
    .CLK(clknet_leaf_163_clock),
    .Q(\stack[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10802_ (.D(_00394_),
    .CLK(clknet_leaf_167_clock),
    .Q(\stack[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10803_ (.D(_00395_),
    .CLK(clknet_leaf_166_clock),
    .Q(\stack[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10804_ (.D(_00396_),
    .CLK(clknet_leaf_171_clock),
    .Q(\stack[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10805_ (.D(_00397_),
    .CLK(clknet_leaf_139_clock),
    .Q(\stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10806_ (.D(_00398_),
    .CLK(clknet_leaf_134_clock),
    .Q(\stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10807_ (.D(_00399_),
    .CLK(clknet_leaf_140_clock),
    .Q(\stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10808_ (.D(_00400_),
    .CLK(clknet_leaf_163_clock),
    .Q(\stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10809_ (.D(_00401_),
    .CLK(clknet_leaf_167_clock),
    .Q(\stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10810_ (.D(_00402_),
    .CLK(clknet_leaf_166_clock),
    .Q(\stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10811_ (.D(_00403_),
    .CLK(clknet_leaf_171_clock),
    .Q(\stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10812_ (.D(_00404_),
    .CLK(clknet_leaf_171_clock),
    .Q(\stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10813_ (.D(_00405_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10814_ (.D(_00406_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10815_ (.D(_00407_),
    .CLK(clknet_leaf_159_clock),
    .Q(\stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10816_ (.D(_00408_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10817_ (.D(_00409_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10818_ (.D(_00410_),
    .CLK(clknet_leaf_168_clock),
    .Q(\stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10819_ (.D(_00411_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10820_ (.D(_00412_),
    .CLK(clknet_leaf_170_clock),
    .Q(\stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10821_ (.D(_00413_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10822_ (.D(_00414_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10823_ (.D(_00415_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10824_ (.D(_00416_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10825_ (.D(_00417_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10826_ (.D(_00418_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10827_ (.D(_00419_),
    .CLK(clknet_leaf_171_clock),
    .Q(\stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10828_ (.D(_00420_),
    .CLK(clknet_leaf_171_clock),
    .Q(\stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10829_ (.D(_00421_),
    .CLK(clknet_leaf_157_clock),
    .Q(\stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10830_ (.D(_00422_),
    .CLK(clknet_leaf_153_clock),
    .Q(\stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10831_ (.D(_00423_),
    .CLK(clknet_leaf_157_clock),
    .Q(\stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10832_ (.D(_00424_),
    .CLK(clknet_leaf_153_clock),
    .Q(\stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10833_ (.D(_00425_),
    .CLK(clknet_leaf_154_clock),
    .Q(\stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10834_ (.D(_00426_),
    .CLK(clknet_leaf_177_clock),
    .Q(\stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10835_ (.D(_00427_),
    .CLK(clknet_leaf_189_clock),
    .Q(\stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10836_ (.D(_00428_),
    .CLK(clknet_leaf_189_clock),
    .Q(\stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10837_ (.D(_00429_),
    .CLK(clknet_leaf_139_clock),
    .Q(\stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10838_ (.D(_00430_),
    .CLK(clknet_leaf_154_clock),
    .Q(\stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10839_ (.D(_00431_),
    .CLK(clknet_leaf_153_clock),
    .Q(\stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10840_ (.D(_00432_),
    .CLK(clknet_leaf_177_clock),
    .Q(\stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10841_ (.D(_00433_),
    .CLK(clknet_leaf_176_clock),
    .Q(\stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10842_ (.D(_00434_),
    .CLK(clknet_leaf_175_clock),
    .Q(\stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10843_ (.D(_00435_),
    .CLK(clknet_leaf_190_clock),
    .Q(\stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10844_ (.D(_00436_),
    .CLK(clknet_leaf_189_clock),
    .Q(\stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10845_ (.D(_00437_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10846_ (.D(_00438_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10847_ (.D(_00439_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10848_ (.D(_00440_),
    .CLK(clknet_leaf_161_clock),
    .Q(\stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10849_ (.D(_00441_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10850_ (.D(_00442_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10851_ (.D(_00443_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10852_ (.D(_00444_),
    .CLK(clknet_leaf_173_clock),
    .Q(\stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10853_ (.D(_00445_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10854_ (.D(_00446_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10855_ (.D(_00447_),
    .CLK(clknet_leaf_160_clock),
    .Q(\stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10856_ (.D(_00448_),
    .CLK(clknet_leaf_162_clock),
    .Q(\stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10857_ (.D(_00449_),
    .CLK(clknet_leaf_168_clock),
    .Q(\stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10858_ (.D(_00450_),
    .CLK(clknet_leaf_168_clock),
    .Q(\stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10859_ (.D(_00451_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10860_ (.D(_00452_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10861_ (.D(_00453_),
    .CLK(clknet_leaf_145_clock),
    .Q(\stack[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10862_ (.D(_00454_),
    .CLK(clknet_leaf_152_clock),
    .Q(\stack[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10863_ (.D(_00455_),
    .CLK(clknet_leaf_144_clock),
    .Q(\stack[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10864_ (.D(_00456_),
    .CLK(clknet_leaf_150_clock),
    .Q(\stack[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10865_ (.D(_00457_),
    .CLK(clknet_leaf_150_clock),
    .Q(\stack[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10866_ (.D(_00458_),
    .CLK(clknet_leaf_183_clock),
    .Q(\stack[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10867_ (.D(_00459_),
    .CLK(clknet_leaf_190_clock),
    .Q(\stack[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10868_ (.D(_00460_),
    .CLK(clknet_leaf_190_clock),
    .Q(\stack[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10869_ (.D(_00461_),
    .CLK(clknet_leaf_140_clock),
    .Q(\stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10870_ (.D(_00462_),
    .CLK(clknet_leaf_152_clock),
    .Q(\stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10871_ (.D(_00463_),
    .CLK(clknet_leaf_145_clock),
    .Q(\stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10872_ (.D(_00464_),
    .CLK(clknet_leaf_152_clock),
    .Q(\stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10873_ (.D(_00465_),
    .CLK(clknet_leaf_149_clock),
    .Q(\stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10874_ (.D(_00466_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10875_ (.D(_00467_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10876_ (.D(_00468_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10877_ (.D(_00469_),
    .CLK(clknet_leaf_144_clock),
    .Q(\stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10878_ (.D(_00470_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10879_ (.D(_00471_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10880_ (.D(_00472_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10881_ (.D(_00473_),
    .CLK(clknet_leaf_179_clock),
    .Q(\stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10882_ (.D(_00474_),
    .CLK(clknet_leaf_183_clock),
    .Q(\stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10883_ (.D(_00475_),
    .CLK(clknet_leaf_193_clock),
    .Q(\stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10884_ (.D(_00476_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10885_ (.D(_00477_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10886_ (.D(_00478_),
    .CLK(clknet_leaf_146_clock),
    .Q(\stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10887_ (.D(_00479_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10888_ (.D(_00480_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10889_ (.D(_00481_),
    .CLK(clknet_leaf_181_clock),
    .Q(\stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10890_ (.D(_00482_),
    .CLK(clknet_leaf_183_clock),
    .Q(\stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10891_ (.D(_00483_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10892_ (.D(_00484_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10893_ (.D(_00485_),
    .CLK(clknet_leaf_146_clock),
    .Q(\stack[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10894_ (.D(_00486_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10895_ (.D(_00487_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10896_ (.D(_00488_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10897_ (.D(_00489_),
    .CLK(clknet_leaf_182_clock),
    .Q(\stack[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10898_ (.D(_00490_),
    .CLK(clknet_leaf_185_clock),
    .Q(\stack[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10899_ (.D(_00491_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10900_ (.D(_00492_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10901_ (.D(_00493_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10902_ (.D(_00494_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10903_ (.D(_00495_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10904_ (.D(_00496_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10905_ (.D(_00497_),
    .CLK(clknet_leaf_181_clock),
    .Q(\stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10906_ (.D(_00498_),
    .CLK(clknet_leaf_185_clock),
    .Q(\stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10907_ (.D(_00499_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10908_ (.D(_00500_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10909_ (.D(_00501_),
    .CLK(clknet_leaf_139_clock),
    .Q(\stack[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10910_ (.D(_00502_),
    .CLK(clknet_leaf_179_clock),
    .Q(\stack[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10911_ (.D(_00503_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10912_ (.D(_00504_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10913_ (.D(_00505_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10914_ (.D(_00506_),
    .CLK(clknet_leaf_184_clock),
    .Q(\stack[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10915_ (.D(_00507_),
    .CLK(clknet_leaf_188_clock),
    .Q(\stack[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10916_ (.D(_00508_),
    .CLK(clknet_leaf_188_clock),
    .Q(\stack[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10917_ (.D(_00509_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10918_ (.D(_00510_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10919_ (.D(_00511_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10920_ (.D(_00512_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10921_ (.D(_00513_),
    .CLK(clknet_leaf_182_clock),
    .Q(\stack[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10922_ (.D(_00514_),
    .CLK(clknet_leaf_185_clock),
    .Q(\stack[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10923_ (.D(_00515_),
    .CLK(clknet_leaf_187_clock),
    .Q(\stack[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10924_ (.D(_00516_),
    .CLK(clknet_leaf_186_clock),
    .Q(\stack[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10925_ (.D(_00517_),
    .CLK(clknet_leaf_34_clock),
    .Q(wb_read_ack));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10926_ (.D(_00518_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10927_ (.D(_00519_),
    .CLK(clknet_leaf_148_clock),
    .Q(\stack[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10928_ (.D(_00520_),
    .CLK(clknet_leaf_147_clock),
    .Q(\stack[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10929_ (.D(_00521_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10930_ (.D(_00522_),
    .CLK(clknet_leaf_182_clock),
    .Q(\stack[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10931_ (.D(_00523_),
    .CLK(clknet_leaf_182_clock),
    .Q(\stack[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10932_ (.D(_00524_),
    .CLK(clknet_leaf_191_clock),
    .Q(\stack[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10933_ (.D(_00525_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10934_ (.D(_00526_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10935_ (.D(_00527_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10936_ (.D(_00528_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10937_ (.D(_00529_),
    .CLK(clknet_leaf_149_clock),
    .Q(\stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10938_ (.D(_00530_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10939_ (.D(_00531_),
    .CLK(clknet_leaf_183_clock),
    .Q(\stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10940_ (.D(_00532_),
    .CLK(clknet_leaf_191_clock),
    .Q(\stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10941_ (.D(_00533_),
    .CLK(clknet_leaf_0_clock),
    .Q(\stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10942_ (.D(_00534_),
    .CLK(clknet_leaf_146_clock),
    .Q(\stack[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10943_ (.D(_00535_),
    .CLK(clknet_leaf_142_clock),
    .Q(\stack[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10944_ (.D(_00536_),
    .CLK(clknet_leaf_142_clock),
    .Q(\stack[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10945_ (.D(_00537_),
    .CLK(clknet_leaf_149_clock),
    .Q(\stack[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10946_ (.D(_00538_),
    .CLK(clknet_leaf_180_clock),
    .Q(\stack[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10947_ (.D(_00539_),
    .CLK(clknet_leaf_182_clock),
    .Q(\stack[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10948_ (.D(_00540_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10949_ (.D(_00541_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10950_ (.D(_00542_),
    .CLK(clknet_leaf_144_clock),
    .Q(\stack[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10951_ (.D(_00543_),
    .CLK(clknet_leaf_143_clock),
    .Q(\stack[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10952_ (.D(_00544_),
    .CLK(clknet_leaf_144_clock),
    .Q(\stack[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10953_ (.D(_00545_),
    .CLK(clknet_leaf_149_clock),
    .Q(\stack[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10954_ (.D(_00546_),
    .CLK(clknet_leaf_179_clock),
    .Q(\stack[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10955_ (.D(_00547_),
    .CLK(clknet_leaf_183_clock),
    .Q(\stack[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10956_ (.D(_00548_),
    .CLK(clknet_leaf_187_clock),
    .Q(\stack[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10957_ (.D(_00549_),
    .CLK(clknet_leaf_187_clock),
    .Q(\stack[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10958_ (.D(_00550_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10959_ (.D(_00551_),
    .CLK(clknet_leaf_142_clock),
    .Q(\stack[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10960_ (.D(_00552_),
    .CLK(clknet_leaf_142_clock),
    .Q(\stack[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10961_ (.D(_00553_),
    .CLK(clknet_leaf_149_clock),
    .Q(\stack[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10962_ (.D(_00554_),
    .CLK(clknet_leaf_179_clock),
    .Q(\stack[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10963_ (.D(_00555_),
    .CLK(clknet_leaf_184_clock),
    .Q(\stack[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10964_ (.D(_00556_),
    .CLK(clknet_leaf_188_clock),
    .Q(\stack[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10965_ (.D(_00557_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10966_ (.D(_00558_),
    .CLK(clknet_leaf_129_clock),
    .Q(net158));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10967_ (.D(_00559_),
    .CLK(clknet_leaf_129_clock),
    .Q(net159));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10968_ (.D(_00560_),
    .CLK(clknet_leaf_43_clock),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10969_ (.D(_00561_),
    .CLK(clknet_4_3_0_clock),
    .Q(net130));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10970_ (.D(_00562_),
    .CLK(clknet_leaf_43_clock),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10971_ (.D(_00563_),
    .CLK(clknet_leaf_43_clock),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10972_ (.D(_00564_),
    .CLK(clknet_4_3_0_clock),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10973_ (.D(_00565_),
    .CLK(clknet_leaf_43_clock),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10974_ (.D(_00566_),
    .CLK(clknet_leaf_42_clock),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10975_ (.D(_00567_),
    .CLK(clknet_leaf_45_clock),
    .Q(net139));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10976_ (.D(_00568_),
    .CLK(clknet_leaf_42_clock),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10977_ (.D(_00569_),
    .CLK(clknet_leaf_44_clock),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10978_ (.D(_00570_),
    .CLK(clknet_leaf_43_clock),
    .Q(net154));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10979_ (.D(_00571_),
    .CLK(clknet_leaf_44_clock),
    .Q(net155));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10980_ (.D(_00572_),
    .CLK(clknet_leaf_44_clock),
    .Q(net156));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10981_ (.D(_00573_),
    .CLK(clknet_leaf_44_clock),
    .Q(net157));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10982_ (.D(_00574_),
    .CLK(clknet_leaf_9_clock),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10983_ (.D(_00575_),
    .CLK(clknet_leaf_9_clock),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10984_ (.D(_00576_),
    .CLK(clknet_4_3_0_clock),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10985_ (.D(_00577_),
    .CLK(clknet_leaf_131_clock),
    .Q(net138));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10986_ (.D(_00578_),
    .CLK(clknet_leaf_9_clock),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10987_ (.D(_00579_),
    .CLK(clknet_leaf_39_clock),
    .Q(\mem.mem_io.past_write ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10988_ (.D(_00580_),
    .CLK(clknet_leaf_13_clock),
    .Q(\exec.out_of_order_exec ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10989_ (.D(_00581_),
    .CLK(clknet_leaf_40_clock),
    .Q(\mem.sram_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10990_ (.D(_00582_),
    .CLK(clknet_leaf_41_clock),
    .Q(\mem.select ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10991_ (.D(_00583_),
    .CLK(clknet_leaf_40_clock),
    .Q(net141));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10992_ (.D(_00584_),
    .CLK(clknet_leaf_13_clock),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10993_ (.D(_00585_),
    .CLK(clknet_leaf_13_clock),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10994_ (.D(_00586_),
    .CLK(clknet_leaf_10_clock),
    .Q(\intr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10995_ (.D(_00587_),
    .CLK(clknet_leaf_7_clock),
    .Q(\intr_enable[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10996_ (.D(_00588_),
    .CLK(clknet_leaf_8_clock),
    .Q(\intr_enable[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10997_ (.D(_00589_),
    .CLK(clknet_leaf_12_clock),
    .Q(edge_interrupts));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10998_ (.D(_00590_),
    .CLK(clknet_leaf_129_clock),
    .Q(\exec.memory_input[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10999_ (.D(_00591_),
    .CLK(clknet_leaf_129_clock),
    .Q(\exec.memory_input[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11000_ (.D(_00592_),
    .CLK(clknet_leaf_128_clock),
    .Q(\exec.memory_input[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11001_ (.D(_00593_),
    .CLK(clknet_leaf_128_clock),
    .Q(\exec.memory_input[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11002_ (.D(_00594_),
    .CLK(clknet_leaf_127_clock),
    .Q(\exec.memory_input[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11003_ (.D(_00595_),
    .CLK(clknet_leaf_128_clock),
    .Q(\exec.memory_input[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11004_ (.D(_00596_),
    .CLK(clknet_leaf_129_clock),
    .Q(\exec.memory_input[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11005_ (.D(_00597_),
    .CLK(clknet_leaf_128_clock),
    .Q(\exec.memory_input[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11006_ (.D(_00598_),
    .CLK(clknet_leaf_12_clock),
    .Q(single_step));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11007_ (.D(_00599_),
    .CLK(clknet_leaf_13_clock),
    .Q(prev_level_interrupt));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11008_ (.D(_00600_),
    .CLK(clknet_leaf_127_clock),
    .Q(\mem.mem_dff.memory_type_data ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11009_ (.D(_00601_),
    .CLK(clknet_leaf_46_clock),
    .Q(\mem.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11010_ (.D(_00602_),
    .CLK(clknet_leaf_45_clock),
    .Q(\mem.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11011_ (.D(_00603_),
    .CLK(clknet_leaf_46_clock),
    .Q(net185));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11012_ (.D(_00604_),
    .CLK(clknet_leaf_127_clock),
    .Q(net186));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11013_ (.D(_00605_),
    .CLK(clknet_4_12_0_clock),
    .Q(net187));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11014_ (.D(_00606_),
    .CLK(clknet_leaf_127_clock),
    .Q(net188));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11015_ (.D(_00607_),
    .CLK(clknet_leaf_127_clock),
    .Q(net189));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11016_ (.D(_00608_),
    .CLK(clknet_leaf_127_clock),
    .Q(net190));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11017_ (.D(_00609_),
    .CLK(clknet_leaf_41_clock),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11018_ (.D(_00610_),
    .CLK(clknet_leaf_17_clock),
    .Q(\cycles_per_ms[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11019_ (.D(_00611_),
    .CLK(clknet_leaf_7_clock),
    .Q(\cycles_per_ms[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11020_ (.D(_00612_),
    .CLK(clknet_leaf_16_clock),
    .Q(\cycles_per_ms[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11021_ (.D(_00613_),
    .CLK(clknet_leaf_16_clock),
    .Q(\cycles_per_ms[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11022_ (.D(_00614_),
    .CLK(clknet_leaf_15_clock),
    .Q(\cycles_per_ms[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11023_ (.D(_00615_),
    .CLK(clknet_leaf_16_clock),
    .Q(\cycles_per_ms[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11024_ (.D(_00616_),
    .CLK(clknet_leaf_17_clock),
    .Q(\cycles_per_ms[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11025_ (.D(_00617_),
    .CLK(clknet_leaf_15_clock),
    .Q(\cycles_per_ms[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11026_ (.D(_00618_),
    .CLK(clknet_leaf_17_clock),
    .Q(\cycles_per_ms[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11027_ (.D(_00619_),
    .CLK(clknet_leaf_17_clock),
    .Q(\cycles_per_ms[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11028_ (.D(_00620_),
    .CLK(clknet_leaf_19_clock),
    .Q(\cycles_per_ms[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11029_ (.D(_00621_),
    .CLK(clknet_leaf_14_clock),
    .Q(\cycles_per_ms[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11030_ (.D(_00622_),
    .CLK(clknet_leaf_20_clock),
    .Q(\cycles_per_ms[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11031_ (.D(_00623_),
    .CLK(clknet_4_8_0_clock),
    .Q(\cycles_per_ms[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11032_ (.D(_00624_),
    .CLK(clknet_leaf_19_clock),
    .Q(\cycles_per_ms[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11033_ (.D(_00625_),
    .CLK(clknet_leaf_19_clock),
    .Q(\cycles_per_ms[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11034_ (.D(_00626_),
    .CLK(clknet_leaf_33_clock),
    .Q(\cycles_per_ms[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11035_ (.D(_00627_),
    .CLK(clknet_leaf_22_clock),
    .Q(\cycles_per_ms[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11036_ (.D(_00628_),
    .CLK(clknet_leaf_32_clock),
    .Q(\cycles_per_ms[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11037_ (.D(_00629_),
    .CLK(clknet_leaf_33_clock),
    .Q(\cycles_per_ms[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11038_ (.D(_00630_),
    .CLK(clknet_leaf_33_clock),
    .Q(\cycles_per_ms[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11039_ (.D(_00631_),
    .CLK(clknet_leaf_33_clock),
    .Q(\cycles_per_ms[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11040_ (.D(_00632_),
    .CLK(clknet_leaf_34_clock),
    .Q(\cycles_per_ms[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11041_ (.D(_00633_),
    .CLK(clknet_leaf_34_clock),
    .Q(\cycles_per_ms[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11042_ (.D(_00634_),
    .CLK(clknet_leaf_17_clock),
    .Q(\delay_cycles[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11043_ (.D(_00635_),
    .CLK(clknet_leaf_26_clock),
    .Q(\delay_cycles[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11044_ (.D(_00636_),
    .CLK(clknet_4_2_0_clock),
    .Q(\delay_cycles[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11045_ (.D(_00637_),
    .CLK(clknet_leaf_26_clock),
    .Q(\delay_cycles[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11046_ (.D(_00638_),
    .CLK(clknet_leaf_26_clock),
    .Q(\delay_cycles[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11047_ (.D(_00639_),
    .CLK(clknet_leaf_26_clock),
    .Q(\delay_cycles[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11048_ (.D(_00640_),
    .CLK(clknet_leaf_26_clock),
    .Q(\delay_cycles[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11049_ (.D(_00641_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11050_ (.D(_00642_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11051_ (.D(_00643_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11052_ (.D(_00644_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11053_ (.D(_00645_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11054_ (.D(_00646_),
    .CLK(clknet_leaf_25_clock),
    .Q(\delay_cycles[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11055_ (.D(_00647_),
    .CLK(clknet_leaf_24_clock),
    .Q(\delay_cycles[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11056_ (.D(_00648_),
    .CLK(clknet_leaf_24_clock),
    .Q(\delay_cycles[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11057_ (.D(_00649_),
    .CLK(clknet_leaf_23_clock),
    .Q(\delay_cycles[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11058_ (.D(_00650_),
    .CLK(clknet_leaf_22_clock),
    .Q(\delay_cycles[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11059_ (.D(_00651_),
    .CLK(clknet_leaf_23_clock),
    .Q(\delay_cycles[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11060_ (.D(_00652_),
    .CLK(clknet_leaf_22_clock),
    .Q(\delay_cycles[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11061_ (.D(_00653_),
    .CLK(clknet_leaf_21_clock),
    .Q(\delay_cycles[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11062_ (.D(_00654_),
    .CLK(clknet_leaf_21_clock),
    .Q(\delay_cycles[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11063_ (.D(_00655_),
    .CLK(clknet_leaf_21_clock),
    .Q(\delay_cycles[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11064_ (.D(_00656_),
    .CLK(clknet_leaf_21_clock),
    .Q(\delay_cycles[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11065_ (.D(_00657_),
    .CLK(clknet_leaf_20_clock),
    .Q(\delay_cycles[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11066_ (.D(_00658_),
    .CLK(clknet_leaf_131_clock),
    .Q(net210));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11067_ (.D(_00659_),
    .CLK(clknet_opt_2_0_clock),
    .Q(net211));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11068_ (.D(_00660_),
    .CLK(clknet_4_0_0_clock),
    .Q(net212));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11069_ (.D(_00661_),
    .CLK(clknet_opt_1_0_clock),
    .Q(net213));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11070_ (.D(_00662_),
    .CLK(clknet_leaf_69_clock),
    .Q(net214));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11071_ (.D(_00663_),
    .CLK(clknet_opt_5_0_clock),
    .Q(net215));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11072_ (.D(_00664_),
    .CLK(clknet_leaf_87_clock),
    .Q(net217));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11073_ (.D(_00665_),
    .CLK(clknet_opt_3_0_clock),
    .Q(net218));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11074_ (.D(_00666_),
    .CLK(clknet_leaf_40_clock),
    .Q(wb_write_ack));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11075_ (.D(_00667_),
    .CLK(clknet_4_9_0_clock),
    .Q(\delay_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11076_ (.D(_00668_),
    .CLK(clknet_leaf_132_clock),
    .Q(\delay_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11077_ (.D(_00669_),
    .CLK(clknet_leaf_132_clock),
    .Q(\delay_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11078_ (.D(_00670_),
    .CLK(clknet_leaf_132_clock),
    .Q(\delay_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11079_ (.D(_00671_),
    .CLK(clknet_leaf_125_clock),
    .Q(\delay_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11080_ (.D(_00672_),
    .CLK(clknet_leaf_125_clock),
    .Q(\delay_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11081_ (.D(_00673_),
    .CLK(clknet_leaf_127_clock),
    .Q(\delay_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11082_ (.D(_00674_),
    .CLK(clknet_leaf_125_clock),
    .Q(\delay_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11083_ (.D(_00675_),
    .CLK(clknet_leaf_40_clock),
    .Q(net161));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11084_ (.D(_00676_),
    .CLK(clknet_leaf_129_clock),
    .Q(net172));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11085_ (.D(_00677_),
    .CLK(clknet_leaf_10_clock),
    .Q(net177));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11086_ (.D(_00678_),
    .CLK(clknet_leaf_10_clock),
    .Q(net178));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11087_ (.D(_00679_),
    .CLK(clknet_leaf_44_clock),
    .Q(net179));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11088_ (.D(_00680_),
    .CLK(clknet_leaf_128_clock),
    .Q(net180));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11089_ (.D(_00681_),
    .CLK(clknet_leaf_15_clock),
    .Q(net181));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11090_ (.D(_00682_),
    .CLK(clknet_leaf_15_clock),
    .Q(net182));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11091_ (.D(_00683_),
    .CLK(clknet_leaf_14_clock),
    .Q(net183));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11092_ (.D(_00684_),
    .CLK(clknet_leaf_14_clock),
    .Q(net184));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11093_ (.D(_00685_),
    .CLK(clknet_leaf_14_clock),
    .Q(net162));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11094_ (.D(_00686_),
    .CLK(clknet_leaf_14_clock),
    .Q(net163));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11095_ (.D(_00687_),
    .CLK(clknet_leaf_6_clock),
    .Q(net164));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11096_ (.D(_00688_),
    .CLK(clknet_leaf_6_clock),
    .Q(net165));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11097_ (.D(_00689_),
    .CLK(clknet_leaf_6_clock),
    .Q(net166));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11098_ (.D(_00690_),
    .CLK(clknet_leaf_14_clock),
    .Q(net167));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11099_ (.D(_00691_),
    .CLK(clknet_leaf_32_clock),
    .Q(net168));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11100_ (.D(_00692_),
    .CLK(clknet_leaf_35_clock),
    .Q(net169));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11101_ (.D(_00693_),
    .CLK(clknet_leaf_33_clock),
    .Q(net170));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11102_ (.D(_00694_),
    .CLK(clknet_leaf_35_clock),
    .Q(net171));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11103_ (.D(_00695_),
    .CLK(clknet_leaf_34_clock),
    .Q(net173));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11104_ (.D(_00696_),
    .CLK(clknet_leaf_34_clock),
    .Q(net174));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11105_ (.D(_00697_),
    .CLK(clknet_leaf_35_clock),
    .Q(net175));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11106_ (.D(_00698_),
    .CLK(clknet_leaf_35_clock),
    .Q(net176));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11107_ (.D(_00699_),
    .CLK(clknet_leaf_8_clock),
    .Q(prev_reg_write));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11108_ (.D(_00700_),
    .CLK(clknet_leaf_144_clock),
    .Q(\stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11109_ (.D(_00701_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11110_ (.D(_00702_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11111_ (.D(_00703_),
    .CLK(clknet_leaf_151_clock),
    .Q(\stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11112_ (.D(_00704_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11113_ (.D(_00705_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11114_ (.D(_00706_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11115_ (.D(_00707_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11116_ (.D(_00708_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11117_ (.D(_00709_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11118_ (.D(_00710_),
    .CLK(clknet_leaf_141_clock),
    .Q(\stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11119_ (.D(_00711_),
    .CLK(clknet_leaf_151_clock),
    .Q(\stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11120_ (.D(_00712_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11121_ (.D(_00713_),
    .CLK(clknet_leaf_178_clock),
    .Q(\stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11122_ (.D(_00714_),
    .CLK(clknet_leaf_189_clock),
    .Q(\stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11123_ (.D(_00715_),
    .CLK(clknet_leaf_192_clock),
    .Q(\stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11124_ (.D(_00716_),
    .CLK(clknet_leaf_158_clock),
    .Q(\stack[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11125_ (.D(_00717_),
    .CLK(clknet_leaf_158_clock),
    .Q(\stack[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11126_ (.D(_00718_),
    .CLK(clknet_leaf_158_clock),
    .Q(\stack[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11127_ (.D(_00719_),
    .CLK(clknet_leaf_156_clock),
    .Q(\stack[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11128_ (.D(_00720_),
    .CLK(clknet_leaf_169_clock),
    .Q(\stack[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11129_ (.D(_00721_),
    .CLK(clknet_leaf_173_clock),
    .Q(\stack[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11130_ (.D(_00722_),
    .CLK(clknet_leaf_173_clock),
    .Q(\stack[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11131_ (.D(_00723_),
    .CLK(clknet_leaf_173_clock),
    .Q(\stack[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11132_ (.D(_00724_),
    .CLK(clknet_leaf_153_clock),
    .Q(\stack[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11133_ (.D(_00725_),
    .CLK(clknet_leaf_152_clock),
    .Q(\stack[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11134_ (.D(_00726_),
    .CLK(clknet_leaf_145_clock),
    .Q(\stack[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11135_ (.D(_00727_),
    .CLK(clknet_leaf_151_clock),
    .Q(\stack[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11136_ (.D(_00728_),
    .CLK(clknet_leaf_179_clock),
    .Q(\stack[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11137_ (.D(_00729_),
    .CLK(clknet_leaf_184_clock),
    .Q(\stack[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11138_ (.D(_00730_),
    .CLK(clknet_leaf_187_clock),
    .Q(\stack[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11139_ (.D(_00731_),
    .CLK(clknet_leaf_193_clock),
    .Q(\stack[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11140_ (.D(_00732_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11141_ (.D(_00733_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11142_ (.D(_00734_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11143_ (.D(_00735_),
    .CLK(clknet_leaf_156_clock),
    .Q(\stack[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11144_ (.D(_00736_),
    .CLK(clknet_leaf_177_clock),
    .Q(\stack[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11145_ (.D(_00737_),
    .CLK(clknet_4_1_0_clock),
    .Q(\stack[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11146_ (.D(_00738_),
    .CLK(clknet_leaf_191_clock),
    .Q(\stack[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11147_ (.D(_00739_),
    .CLK(clknet_leaf_191_clock),
    .Q(\stack[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11148_ (.D(_00740_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11149_ (.D(_00741_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11150_ (.D(_00742_),
    .CLK(clknet_leaf_138_clock),
    .Q(\stack[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11151_ (.D(_00743_),
    .CLK(clknet_4_7_0_clock),
    .Q(\stack[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11152_ (.D(_00744_),
    .CLK(clknet_leaf_176_clock),
    .Q(\stack[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11153_ (.D(_00745_),
    .CLK(clknet_leaf_175_clock),
    .Q(\stack[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11154_ (.D(_00746_),
    .CLK(clknet_leaf_191_clock),
    .Q(\stack[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11155_ (.D(_00747_),
    .CLK(clknet_leaf_190_clock),
    .Q(\stack[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11156_ (.D(_00748_),
    .CLK(clknet_leaf_133_clock),
    .Q(\stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11157_ (.D(_00749_),
    .CLK(clknet_leaf_133_clock),
    .Q(\stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11158_ (.D(_00750_),
    .CLK(clknet_leaf_133_clock),
    .Q(\stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11159_ (.D(_00751_),
    .CLK(clknet_leaf_168_clock),
    .Q(\stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11160_ (.D(_00752_),
    .CLK(clknet_leaf_167_clock),
    .Q(\stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11161_ (.D(_00753_),
    .CLK(clknet_leaf_166_clock),
    .Q(\stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11162_ (.D(_00754_),
    .CLK(clknet_leaf_5_clock),
    .Q(\stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11163_ (.D(_00755_),
    .CLK(clknet_leaf_5_clock),
    .Q(\stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11175_ (.I(clknet_opt_4_1_clock),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11176_ (.I(net249),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11177_ (.I(net247),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11178_ (.I(net244),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11179_ (.I(net242),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11180_ (.I(net240),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11181_ (.I(net237),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11182_ (.I(net235),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11183_ (.I(net233),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11184_ (.I(net250),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11185_ (.I(net247),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11186_ (.I(net245),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11187_ (.I(net243),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11188_ (.I(net241),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11189_ (.I(net237),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11190_ (.I(net235),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11191_ (.I(net234),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11192_ (.I(net251),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11193_ (.I(net247),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11194_ (.I(net246),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11195_ (.I(net242),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11196_ (.I(net241),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11197_ (.I(net238),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11198_ (.I(net236),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11199_ (.I(net233),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11200_ (.I(net110),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11201_ (.I(net193),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input1 (.I(i_la_addr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(i_la_addr[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(i_la_addr[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(i_la_addr[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(i_la_addr[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(i_la_addr[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(i_la_addr[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(i_la_data[0]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(i_la_data[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(i_la_data[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(i_la_data[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(i_la_data[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(i_la_data[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(i_la_data[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(i_la_data[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input16 (.I(i_la_wb_disable),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(i_la_write),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input18 (.I(i_wb_addr[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(i_wb_addr[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(i_wb_addr[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input21 (.I(i_wb_addr[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input22 (.I(i_wb_addr[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input23 (.I(i_wb_addr[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(i_wb_addr[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(i_wb_addr[16]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(i_wb_addr[17]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(i_wb_addr[18]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(i_wb_addr[19]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(i_wb_addr[1]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(i_wb_addr[20]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input31 (.I(i_wb_addr[21]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(i_wb_addr[22]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(i_wb_addr[23]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(i_wb_addr[2]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(i_wb_addr[3]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(i_wb_addr[4]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input37 (.I(i_wb_addr[5]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(i_wb_addr[6]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input39 (.I(i_wb_addr[7]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input40 (.I(i_wb_addr[8]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input41 (.I(i_wb_addr[9]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(i_wb_cyc),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(i_wb_data[0]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input44 (.I(i_wb_data[10]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input45 (.I(i_wb_data[11]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input46 (.I(i_wb_data[12]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input47 (.I(i_wb_data[13]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input48 (.I(i_wb_data[14]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input49 (.I(i_wb_data[15]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input50 (.I(i_wb_data[16]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(i_wb_data[17]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input52 (.I(i_wb_data[18]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(i_wb_data[19]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input54 (.I(i_wb_data[1]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input55 (.I(i_wb_data[20]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input56 (.I(i_wb_data[21]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input57 (.I(i_wb_data[22]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(i_wb_data[23]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input59 (.I(i_wb_data[2]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(i_wb_data[3]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input61 (.I(i_wb_data[4]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input62 (.I(i_wb_data[5]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input63 (.I(i_wb_data[6]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input64 (.I(i_wb_data[7]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(i_wb_data[8]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(i_wb_data[9]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(i_wb_stb),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input68 (.I(i_wb_we),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(io_in[0]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(io_in[1]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input71 (.I(io_in[2]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(io_in[3]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input73 (.I(io_in[4]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(io_in[5]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input75 (.I(io_in[6]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input76 (.I(io_in[7]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input77 (.I(rambus_wb_ack_i),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input78 (.I(rambus_wb_dat_i[0]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input79 (.I(rambus_wb_dat_i[10]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(rambus_wb_dat_i[11]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input81 (.I(rambus_wb_dat_i[12]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input82 (.I(rambus_wb_dat_i[13]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input83 (.I(rambus_wb_dat_i[14]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input84 (.I(rambus_wb_dat_i[15]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input85 (.I(rambus_wb_dat_i[16]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input86 (.I(rambus_wb_dat_i[17]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input87 (.I(rambus_wb_dat_i[18]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input88 (.I(rambus_wb_dat_i[19]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input89 (.I(rambus_wb_dat_i[1]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(rambus_wb_dat_i[20]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input91 (.I(rambus_wb_dat_i[21]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input92 (.I(rambus_wb_dat_i[22]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input93 (.I(rambus_wb_dat_i[23]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input94 (.I(rambus_wb_dat_i[24]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(rambus_wb_dat_i[25]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input96 (.I(rambus_wb_dat_i[26]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input97 (.I(rambus_wb_dat_i[27]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input98 (.I(rambus_wb_dat_i[28]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(rambus_wb_dat_i[29]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input100 (.I(rambus_wb_dat_i[2]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(rambus_wb_dat_i[30]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(rambus_wb_dat_i[31]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input103 (.I(rambus_wb_dat_i[3]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input104 (.I(rambus_wb_dat_i[4]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input105 (.I(rambus_wb_dat_i[5]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input106 (.I(rambus_wb_dat_i[6]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input107 (.I(rambus_wb_dat_i[7]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input108 (.I(rambus_wb_dat_i[8]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input109 (.I(rambus_wb_dat_i[9]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input110 (.I(reset),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output111 (.I(net111),
    .Z(interrupt));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output112 (.I(net112),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output113 (.I(net113),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output114 (.I(net114),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output115 (.I(net115),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output116 (.I(net116),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output117 (.I(net117),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output118 (.I(net118),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output119 (.I(net119),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output120 (.I(net120),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output121 (.I(net121),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output122 (.I(net122),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output123 (.I(net123),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output124 (.I(net124),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output125 (.I(net125),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output126 (.I(net126),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output131 (.I(net131),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output132 (.I(net132),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net256),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net258),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(o_wb_ack));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(o_wb_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(o_wb_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(o_wb_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(o_wb_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(o_wb_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(o_wb_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(o_wb_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(o_wb_data[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(o_wb_data[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(o_wb_data[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(o_wb_data[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(o_wb_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(o_wb_data[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(o_wb_data[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(o_wb_data[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(o_wb_data[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(o_wb_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(o_wb_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(o_wb_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(o_wb_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(o_wb_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(o_wb_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(o_wb_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(o_wb_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(rambus_wb_addr_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net254),
    .Z(rambus_wb_addr_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(rambus_wb_addr_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(rambus_wb_addr_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(rambus_wb_addr_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(rambus_wb_addr_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(rambus_wb_addr_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 output192 (.I(net192),
    .Z(rambus_wb_clk_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output193 (.I(net193),
    .Z(rambus_wb_cyc_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output194 (.I(net194),
    .Z(rambus_wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output195 (.I(net195),
    .Z(rambus_wb_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output196 (.I(net196),
    .Z(rambus_wb_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output197 (.I(net197),
    .Z(rambus_wb_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output198 (.I(net198),
    .Z(rambus_wb_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output199 (.I(net199),
    .Z(rambus_wb_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output200 (.I(net200),
    .Z(rambus_wb_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output201 (.I(net201),
    .Z(rambus_wb_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output202 (.I(net202),
    .Z(rambus_wb_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output203 (.I(net203),
    .Z(rambus_wb_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output204 (.I(net204),
    .Z(rambus_wb_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output205 (.I(net205),
    .Z(rambus_wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output206 (.I(net206),
    .Z(rambus_wb_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output207 (.I(net207),
    .Z(rambus_wb_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output208 (.I(net208),
    .Z(rambus_wb_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output209 (.I(net209),
    .Z(rambus_wb_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output210 (.I(net252),
    .Z(rambus_wb_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output211 (.I(net248),
    .Z(rambus_wb_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output212 (.I(net246),
    .Z(rambus_wb_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output213 (.I(net243),
    .Z(rambus_wb_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output214 (.I(net240),
    .Z(rambus_wb_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output215 (.I(net239),
    .Z(rambus_wb_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output216 (.I(net216),
    .Z(rambus_wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output217 (.I(net236),
    .Z(rambus_wb_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output218 (.I(net234),
    .Z(rambus_wb_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output219 (.I(net219),
    .Z(rambus_wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output220 (.I(net220),
    .Z(rambus_wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output221 (.I(net221),
    .Z(rambus_wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output222 (.I(net222),
    .Z(rambus_wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output223 (.I(net223),
    .Z(rambus_wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output224 (.I(net224),
    .Z(rambus_wb_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output225 (.I(net225),
    .Z(rambus_wb_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output226 (.I(net226),
    .Z(rambus_wb_rst_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output227 (.I(net227),
    .Z(rambus_wb_sel_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output228 (.I(net228),
    .Z(rambus_wb_sel_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output229 (.I(net229),
    .Z(rambus_wb_sel_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output230 (.I(net230),
    .Z(rambus_wb_sel_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output231 (.I(net231),
    .Z(rambus_wb_stb_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output232 (.I(net253),
    .Z(rambus_wb_we_o));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout233 (.I(net234),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout234 (.I(net218),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout235 (.I(net217),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout236 (.I(net217),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout237 (.I(net239),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout238 (.I(net239),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout239 (.I(net215),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout240 (.I(net241),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout241 (.I(net214),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout242 (.I(net243),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout243 (.I(net213),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout244 (.I(net245),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout245 (.I(net246),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout246 (.I(net212),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout247 (.I(net248),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout248 (.I(net211),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout249 (.I(net250),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout250 (.I(net251),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout251 (.I(net252),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout252 (.I(net210),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout253 (.I(net232),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout254 (.I(net186),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout255 (.I(net185),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout256 (.I(net142),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout257 (.I(net150),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout258 (.I(net159),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel spell_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_6_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_7_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_10_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_12_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_15_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_20_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_21_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_22_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_23_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_24_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_32_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clock (.I(clknet_4_8_0_clock),
    .Z(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_44_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_45_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_46_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_47_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_58_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_65_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_leaf_66_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_71_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_74_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clock (.I(clknet_4_14_0_clock),
    .Z(clknet_leaf_77_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_78_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_80_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_84_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_88_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_89_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_91_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_93_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clock (.I(clknet_4_15_0_clock),
    .Z(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_98_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_107_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_109_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_clock (.I(clknet_4_13_0_clock),
    .Z(clknet_leaf_111_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_114_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_118_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_119_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_124_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clock (.I(clknet_4_9_0_clock),
    .Z(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_131_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clock (.I(clknet_opt_6_0_clock),
    .Z(clknet_leaf_132_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_133_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_134_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_140_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_142_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_144_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_145_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_146_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_150_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_151_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_152_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_clock (.I(clknet_4_5_0_clock),
    .Z(clknet_leaf_154_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_156_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_157_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_clock (.I(clknet_4_6_0_clock),
    .Z(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_166_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_171_clock (.I(clknet_4_3_0_clock),
    .Z(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_175_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_176_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_176_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_177_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_181_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_182_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_182_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_183_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_184_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_184_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_clock (.I(clknet_4_4_0_clock),
    .Z(clknet_leaf_185_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_188_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_189_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_clock (.I(clknet_4_1_0_clock),
    .Z(clknet_leaf_193_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clock (.I(clock),
    .Z(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_0_0_clock (.I(clknet_0_clock),
    .Z(clknet_2_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_1_0_clock (.I(clknet_0_clock),
    .Z(clknet_2_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_2_0_clock (.I(clknet_0_clock),
    .Z(clknet_2_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_3_0_clock (.I(clknet_0_clock),
    .Z(clknet_2_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_clock (.I(clknet_2_0_0_clock),
    .Z(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_clock (.I(clknet_2_0_0_clock),
    .Z(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_clock (.I(clknet_2_1_0_clock),
    .Z(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_clock (.I(clknet_2_1_0_clock),
    .Z(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_clock (.I(clknet_2_2_0_clock),
    .Z(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_clock (.I(clknet_2_2_0_clock),
    .Z(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_clock (.I(clknet_2_3_0_clock),
    .Z(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_clock (.I(clknet_2_3_0_clock),
    .Z(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_clock (.I(clknet_3_0_0_clock),
    .Z(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_clock (.I(clknet_3_0_0_clock),
    .Z(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_clock (.I(clknet_3_1_0_clock),
    .Z(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_clock (.I(clknet_3_1_0_clock),
    .Z(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_clock (.I(clknet_3_2_0_clock),
    .Z(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_clock (.I(clknet_3_2_0_clock),
    .Z(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_clock (.I(clknet_3_3_0_clock),
    .Z(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_clock (.I(clknet_3_3_0_clock),
    .Z(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_clock (.I(clknet_3_4_0_clock),
    .Z(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_clock (.I(clknet_3_4_0_clock),
    .Z(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_clock (.I(clknet_3_5_0_clock),
    .Z(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_clock (.I(clknet_3_5_0_clock),
    .Z(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_clock (.I(clknet_3_6_0_clock),
    .Z(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_clock (.I(clknet_3_6_0_clock),
    .Z(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_clock (.I(clknet_3_7_0_clock),
    .Z(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_clock (.I(clknet_3_7_0_clock),
    .Z(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_clock (.I(clknet_4_0_0_clock),
    .Z(clknet_opt_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_clock (.I(clknet_4_2_0_clock),
    .Z(clknet_opt_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_clock (.I(clknet_4_7_0_clock),
    .Z(clknet_opt_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_0_clock (.I(clknet_4_10_0_clock),
    .Z(clknet_opt_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_1_clock (.I(clknet_opt_4_0_clock),
    .Z(clknet_opt_4_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_5_0_clock (.I(clknet_4_11_0_clock),
    .Z(clknet_opt_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_6_0_clock (.I(clknet_4_12_0_clock),
    .Z(clknet_opt_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__D (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__D (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__D (.I(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__D (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__D (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__D (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__D (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__D (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__D (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__D (.I(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__D (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__D (.I(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__D (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__D (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__D (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__D (.I(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A1 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A1 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A2 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05210__I (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__I (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05212__I (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05459__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05337__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05301__I (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05265__I (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__A3 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05214__I (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05272__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05215__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__S (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__S (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__S (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__A2 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__I (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05221__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05221__A3 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A2 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__A2 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__I (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__B (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__I (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__A2 (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__B2 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__B2 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05224__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05319__B (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__I (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05398__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05283__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05282__B (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A2 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__A2 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05228__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05346__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05242__I (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__S0 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05388__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05236__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__S (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__S (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__S (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__I (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__S (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__S (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__S0 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__S0 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__S1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__S1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__S1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__S1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__S1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__I (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__I (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05262__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__S0 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__S0 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__S (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05246__I (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__S (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__I (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__S0 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__S0 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__S1 (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__I (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__I (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__I (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__B2 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A1 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__S1 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__S1 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__A2 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__S (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__S (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05289__I (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__I (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__S (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__S0 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__S0 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__S0 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__S (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__S (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__S0 (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__I (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__S (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__S0 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S0 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__S0 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__S1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__S1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__S1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__S1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__A2 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__S0 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__S (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__I (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S0 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__S1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__S1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__S1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__A3 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__A2 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__S0 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__S0 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05281__A2 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05284__I (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A1 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A1 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__I (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05285__I (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__B2 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__B2 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__I (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__S (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S0 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__S0 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__S0 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__B2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__C (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__S1 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__S1 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__S1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__S1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__A2 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__A1 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05427__I (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__C (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__B (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__S0 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__S0 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__S0 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__I (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__S (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__S (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__S0 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__S0 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__A2 (.I(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05306__A3 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__A2 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05318__A2 (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__S0 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__S0 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__S (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__S0 (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__S1 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__S1 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__S1 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__S1 (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__A3 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A2 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__I (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__B2 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05323__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__B2 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__B2 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__I (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__B (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__B (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__C (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__A1 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__S (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__I (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05374__I (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__I (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__S (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__S (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__S0 (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__S0 (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__S1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__I (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__S1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__S1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__I0 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__I1 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__I (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__I (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__I (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__S (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__A1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__A1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__A1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__A1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__S1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__S1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__S1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05338__I (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__B2 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__S1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__S1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05354__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__B (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A1 (.I(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__S (.I(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__I (.I(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__S (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__S (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__S0 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__S0 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__S1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__I (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__S1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__S1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05354__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__B (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__C (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05368__I (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__C (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__A2 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__B (.I(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A3 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__I (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__I (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__B2 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A1 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A1 (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__I (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__B2 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__I (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__I (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05540__I (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__B (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__C (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05397__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__A1 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__A1 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__A1 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05384__A1 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__A1 (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__I (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__I (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__I (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__I (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__A1 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A1 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__A1 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__I (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__I (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__S (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A2 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__A1 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__A1 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__I (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__B2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__S1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__B2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__A2 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__A1 (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__I (.I(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05544__I (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__I (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__I (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__A1 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05499__I (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__B1 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__A1 (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__I (.I(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__I (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__A1 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__B1 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05384__A3 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__C (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A1 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__S (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__I (.I(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__I (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__A1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__S (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__S0 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__S (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__B1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__B (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__B2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05394__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05416__I (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05394__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05514__I (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__B1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__B2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__I (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05571__A1 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05449__A1 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05406__A1 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S0 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S0 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__S0 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__S1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__B (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__A2 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05442__I (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__B1 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__I (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__I (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__B1 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__B1 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__A2 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__C (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05478__I (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__C (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__B (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__B2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__B2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__I (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__I (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__S1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__S1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__B2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__C (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__A1 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__S0 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__S0 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__S0 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__I (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__S1 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__S1 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__S1 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__C (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__I (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__B (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05503__I (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__C (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__B (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__A2 (.I(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05522__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__A1 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__B2 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A4 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__I (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__B2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__B2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05432__I (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__I (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05435__A1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__B2 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__A2 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05491__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A1 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__A1 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A1 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05461__I (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__A1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05534__I (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05492__I (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__A1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__S (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__S (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__S (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__I (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05535__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__B2 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A1 (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__I (.I(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__B2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__B2 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__I (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05564__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__S0 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__S0 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05480__I (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__S0 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A1 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__S0 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__S1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__B2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__B2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__S1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A2 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__B1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__B1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05485__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A1 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__A1 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__A1 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__A1 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__C (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__C (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05533__C (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A1 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__I (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05554__I (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__A1 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__A1 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__B2 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__I (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__B2 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__B2 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__I (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__A2 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__B1 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__A2 (.I(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__A2 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05531__I (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__A1 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__A2 (.I(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__C (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__C (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__C (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__C (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__C (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05551__C (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__C (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__A2 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05511__B (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__I (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__A2 (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05537__A1 (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__A2 (.I(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__B2 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__B (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__B1 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__B2 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A2 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__I (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__I (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__B2 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__B2 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A1 (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__I (.I(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__B1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__B1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05533__A1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__B1 (.I(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__B2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__B2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__B2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__B2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__B1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__I (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__I (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__B2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__B2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A1 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__B (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__I (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__C (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__B (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05592__I (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05567__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__B1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__B1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__B (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__I (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A3 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__B1 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__B1 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A2 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__I (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__S0 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__B2 (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A1 (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__S1 (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__B2 (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05573__I (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A2 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A1 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__B2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__I (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A1 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05575__I (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__I (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__I (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__I (.I(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A1 (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__B2 (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__B (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05619__A1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__A1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__C (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__A1 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A1 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__B2 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__B2 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__B2 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__B2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A1 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__A1 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__A1 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__C (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05612__C (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__C (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__C (.I(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__B (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__C (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__A1 (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__B2 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__B2 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__B2 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__I (.I(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05621__I (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__B2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__B2 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__I (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A2 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__A1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A3 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A2 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A3 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A2 (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__B (.I(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__I (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__I (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__B (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__I (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A1 (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A1 (.I(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05661__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__I (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__A1 (.I(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__A1 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A2 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__A2 (.I(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__A2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__A1 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05702__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__I (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A3 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__C (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__I (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A1 (.I(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A1 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__A2 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__A2 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A2 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__I (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05706__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__B (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05682__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A1 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__A2 (.I(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A2 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__A1 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__I (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A3 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__I (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__B (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__B (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__A1 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__B (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A2 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A1 (.I(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A4 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A1 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A2 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05702__B1 (.I(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A2 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__I (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__A3 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__B2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A3 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__A2 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05854__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__A1 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__I (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A1 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__I (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__A1 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__A1 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__S (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__S0 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A2 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__I (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__I (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A1 (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__I (.I(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__B (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A2 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__I (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__A2 (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__I (.I(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A1 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__B2 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__B2 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__B (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__C (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__C (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__A1 (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__B (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__I (.I(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__C (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__I (.I(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__A1 (.I(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__I (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__I (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__B2 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__I (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__B2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__B2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__B2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__B2 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__B2 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__I (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__I (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A1 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A1 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__B2 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__A2 (.I(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A2 (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__B2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__B (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__B2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__I (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__A2 (.I(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__B1 (.I(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__B (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__I (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__I (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__C (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__C (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__I (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__C (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__C (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__C (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__C (.I(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__C (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__C (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__B1 (.I(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__I1 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__B2 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__B (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__S (.I(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__A1 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__A2 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__S (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__S (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__S (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__A1 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__S (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__S0 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__S (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__A2 (.I(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__B1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__B2 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__B2 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__B1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A2 (.I(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__C (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__B (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__C (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__S (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__S (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__S (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__S (.I(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__B1 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__B2 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A1 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__B2 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__B1 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__S (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__S (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__S (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__S (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__S0 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__S (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__S (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__S (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__B1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__S (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__S (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__S (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__S (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__B1 (.I(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A1 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__B1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__A2 (.I(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__B1 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__B2 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__S (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__S (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__S (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__S (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__B2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__B2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__B2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__B2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A2 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A1 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__S (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__S (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__S (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__S (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A1 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__B2 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__B2 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A3 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A1 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__S (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__S (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__S (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__S (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A2 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__S (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__S (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__S (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__S (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__B1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__B2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__B2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__B2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__B2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A2 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__B2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__S (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__S (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__S (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__S (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__B1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__B2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__B2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__B2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__B2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__C (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__C (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__C (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__C (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__B (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__B (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__B (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__B (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__A3 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__S (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__S (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__S (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__S (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__B2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__B2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__B2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__B2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__B2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__B (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__B2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__B2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__S (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__S (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__S (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__S0 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A2 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__S (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__S (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__S (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__S (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__A3 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__A3 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A1 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__S (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__S (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__S (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__S (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A2 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__B (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__S (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__S (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__S (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__S (.I(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__B1 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__B2 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__C (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__C (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__C (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__B1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A4 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__A2 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A3 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A2 (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A2 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A2 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A3 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__A2 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__B1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A2 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A3 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A3 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__B (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__I (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__B2 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A2 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A2 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A2 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__B (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__B1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A1 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A2 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A2 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A2 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__B1 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A3 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A3 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__B (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A3 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A3 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__I (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__S (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__I (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A2 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__B (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A2 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A1 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A1 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A2 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__C (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A2 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A2 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__B (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__I (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__B2 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__S (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__S (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__S (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A1 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A2 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A2 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A1 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__B (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A2 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A2 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__I (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__I (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__S (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__I (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__I (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__I (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A3 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A3 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A3 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A4 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A4 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__B2 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__B2 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__I (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A2 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A2 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A2 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A3 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A2 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A2 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A2 (.I(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__B (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__A1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__B (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__B2 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__B2 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__B2 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__B2 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A2 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A2 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__I (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__I (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__I (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__B2 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__I (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__B1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A1 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__I (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__I (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__I (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A2 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A3 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A3 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__B1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__I (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__I (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__B1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__I (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__I (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__B1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__I (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__B2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A1 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__B2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__B (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A1 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A2 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__B (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__B (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__B (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__I (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__B (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__B1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__B1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__I (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__I (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__I (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__I (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A2 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__B2 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__B1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__I (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__I (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__B1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__I (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A3 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__B2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__B (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__B1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__I (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__I (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__I (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A1 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__B1 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__I (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__I (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A3 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__I (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__I (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__B (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A2 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__B1 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__I (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__I (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__B2 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__I (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__C (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__B2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A2 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A2 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A2 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__I (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__I (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__I (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__I (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__I (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__I (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__I (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__I (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A1 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__B (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__B (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__I (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__I (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__I (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__B (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__B (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__I (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__I (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__I (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__C (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__C (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__C (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__I (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__I (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__I (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A1 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A1 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__I (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A1 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__C (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__C (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__C (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A2 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__I (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__I (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__I (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__I (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__B (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__B (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__B (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__I (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__I (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__I (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__I (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A1 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A1 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__B (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__B (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__B (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__B (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A3 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A3 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A2 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A1 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A3 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A1 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A3 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A3 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A2 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__I (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__I (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__I (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A2 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__I (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__C (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__I (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__B1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__B1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__B1 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A2 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A4 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A2 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A2 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__I (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__I (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__I (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__I (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__I (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__I (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A1 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A1 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A1 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__B (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__B (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__B (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__B (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A3 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A1 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A3 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A2 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__B1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__I (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A3 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A3 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__I (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__I (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__I (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__B (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__B (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__B (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__B (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__B (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__B (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__B (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__B (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__B (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__B (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__B (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__B (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__B (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A1 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A1 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A1 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A1 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__B (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__B (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__B (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__B (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__I (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__I (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__I (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__I (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__I (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__I (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__B (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__B (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__B (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__B (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__B (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__B (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__B (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__B (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__B (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__I (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__I (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__B (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__B (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__B (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__B (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__B (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__B (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A3 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__I (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__I (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A2 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A1 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__B (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__B (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__B (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__B (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__B1 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__I (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A2 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__B1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__A2 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A2 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A2 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__B (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__B (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__B (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__B (.I(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__B1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__B1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__I (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__B1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__B1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__B1 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__I (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__B1 (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__B1 (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__B1 (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__B (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A3 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__B1 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__I (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A1 (.I(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__B (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__B (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__B (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__B (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__I (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A1 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__B (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__B (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__B (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__B (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__I (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__I (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__I (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__I (.I(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A2 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__B (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__B (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__B (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__B (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__B (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__B1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A3 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__B1 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__B1 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__B1 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__B (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__B1 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__B1 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A4 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A2 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A2 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A1 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__B (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__B (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__B (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__B (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__B1 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__I (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__I (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__I (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__B1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__I (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__C2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__C2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__C2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__B (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__B (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__B (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__B (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A1 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__B (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A1 (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A1 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A1 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__B (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__B (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__B (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__B (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A1 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__B1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__I (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__I (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__I (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__I (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A2 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__I (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__B (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__B (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__B (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__B (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__C2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__I (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__I (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__B1 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__B1 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__B1 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__I (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__I (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__I (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__I (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__B1 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__B (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__B (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__B (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__B (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A1 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A1 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A1 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__B1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__B1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__B1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__I (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__I (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__I (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__I (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__B (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__B (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__B (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__B (.I(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__B1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__I (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__B (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__B (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__B (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__B (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__B1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__C2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__B1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__B (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__B (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__B (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__B (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__B (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__B (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__B (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__B (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__B (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__B (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__B (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__B (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A1 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__I (.I(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__I (.I(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__I (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__I (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A1 (.I(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__B (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__B (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__B (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__B (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__B1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__B1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A2 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__I (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A2 (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__I (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__B (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__B (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__B (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__B (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A2 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__I (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__I (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__B (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__B (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__B (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__B (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__B1 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__B2 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__B2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__B (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__B (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__B (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__B2 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__B2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__B (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__B (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__B (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__B (.I(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A2 (.I(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__I (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__I (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__B2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__B2 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__B (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__B (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__B (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__B (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__B2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A1 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__B2 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__B1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__I (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__I (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__B (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__B (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__B (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__B (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__B (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__B (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__B (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__B (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__I (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__I (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__I (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__B (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__B (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__B (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__B (.I(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__B (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__I (.I(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__B (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__B (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__B (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__B (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__B (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__B (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__B (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__B (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A4 (.I(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A4 (.I(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A4 (.I(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A4 (.I(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__I (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A3 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A3 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A3 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A1 (.I(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A3 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__I (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__B1 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__B1 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__B1 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__I (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__B1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__I (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__I (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__I (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A1 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__B1 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A4 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__I (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A4 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__I (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__I (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__I (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A3 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__I (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__I (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__I (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__I (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__I (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__I (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__I (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__C (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__C (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__C (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__B1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__B1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__B1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__B (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__I (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__I (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__I (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I (.I(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__B (.I(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__B (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__I (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__I (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__B1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__C2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__C2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__C2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__B1 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A3 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A3 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__C (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A3 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A4 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__I (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__C (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__I (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__S (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__S (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__S (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__S (.I(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A3 (.I(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A3 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A2 (.I(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__B1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__B1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__B1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__B1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__B1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A4 (.I(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A1 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__B1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__C2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A3 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A4 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__B (.I(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__C (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__C (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__C (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__C (.I(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A3 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__C (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__B1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__B1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__B1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__B1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A3 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__B1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A4 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A4 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A3 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__C (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__C (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B1 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__B1 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__B1 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__B1 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A4 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__B1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A1 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A4 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A3 (.I(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__B2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A3 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__C (.I(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A3 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B1 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A3 (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A3 (.I(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A4 (.I(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__C (.I(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A4 (.I(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B2 (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A1 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A2 (.I(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__C (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__I1 (.I(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__S (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__S (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__S (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__S (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__C (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A2 (.I(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A3 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A4 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__B1 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A3 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A4 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A3 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A4 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__B2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__C (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__I1 (.I(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__C (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A4 (.I(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__B1 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A4 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A3 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__B2 (.I(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A3 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__C (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__I1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__C (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A3 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A4 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__B1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A3 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A4 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A3 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A4 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__B2 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A1 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__C (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__I (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__C (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__C (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__C (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A4 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A3 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A4 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__B (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__I (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__I (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__I (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__I (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__I (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__I (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__I (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A1 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__I (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__I (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A1 (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__B (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__I (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__I (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A1 (.I(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A2 (.I(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__C (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A2 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__C (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__B (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__C (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__C (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__I (.I(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__I (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__I (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__I (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__I (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A2 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A3 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__I (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__B1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__B1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__B1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__B1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A4 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__I (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A2 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A2 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A4 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A4 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A4 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A4 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A2 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A3 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__I (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__I (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__B1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__B1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__B1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A4 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A4 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__I (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A1 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A1 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__B (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A2 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A3 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__I (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A4 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A4 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A4 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A4 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__B1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__I (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__I (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__I (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__I (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__I (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__I (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__I (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__I (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__I (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__I (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__B2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__B2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__I (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A2 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__I (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__I (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A3 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A2 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A2 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A2 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A2 (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__B1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__B1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__B1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__B1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__B1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__B1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__B1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__B1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__I (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A3 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__I (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__B1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__B1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__B1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__B1 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__B1 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B1 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__B1 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A2 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A3 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__B1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__B1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__B1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__B1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__I (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A3 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A3 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A3 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A3 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__I (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A1 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__B1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__B1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__B1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__I (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__I (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__I (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__B2 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__I (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__I (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__I (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__B2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__B2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__B2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__B2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A2 (.I(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__B1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__B1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__B2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__B2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__B2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__B2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__I (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__B1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__B1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__B1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__B1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__B1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A1 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__I (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__B1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__B1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__B1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__B1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__B1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__B1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A2 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__B1 (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__I (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__B1 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__I (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A3 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A3 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A3 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A3 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A4 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A4 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A4 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A4 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__I (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A3 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B1 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__B1 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__B1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__B1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__B1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__B1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__B1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A2 (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__I (.I(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A3 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__B1 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__B1 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__B1 (.I(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__B1 (.I(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__B1 (.I(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__B1 (.I(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__B2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__B2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__B2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A2 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A2 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__I (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A3 (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A3 (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A3 (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A3 (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A2 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A3 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__B1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__B1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A1 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A2 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A3 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__I (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__I (.I(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A2 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__I (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__B1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__B1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__B1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__B1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__B1 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__B1 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__B1 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__B1 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A1 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__I (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__B1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A3 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__B1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__I (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__B1 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A3 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__B1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__B1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__B1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__B1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__B1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__B1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__I (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__I (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__B1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__B1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__B1 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__B1 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__B1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__B2 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__B2 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__B2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__B2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__B1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__I (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A2 (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A2 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A3 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__B1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__B1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__B1 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__B1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A1 (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__C (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__C (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__I (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A3 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__I (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__I (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__I (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A2 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__B1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__B1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__B1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__I (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__B1 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A3 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__B1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__B1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__B1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A2 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A2 (.I(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__B2 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__B2 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__B2 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__B2 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__I (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A1 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A1 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__B1 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__B1 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B1 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__B1 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__I (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__B1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__B1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__B1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__I (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__B1 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A2 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__B1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__B1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__B1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__B1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A2 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A2 (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A1 (.I(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A1 (.I(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__B1 (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__I (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__I (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__A2 (.I(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A2 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__B1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__B1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A1 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__B1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__B1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__B1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__B1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A3 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__I (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__I (.I(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A2 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A2 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A2 (.I(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__B1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__B1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__B1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__B1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__B1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__B1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__B1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A3 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A4 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A3 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A3 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A2 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A3 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__B (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__C (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__I (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__B (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__I (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__C (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A1 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__I (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__I1 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A2 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__B (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__B2 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__C (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__C (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A1 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A1 (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__I1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__I (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__I (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__I (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__C (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__C (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__C (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__C (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__B1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__B1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__B1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__I1 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__C (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__C (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__C (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__C (.I(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A3 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A3 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__B (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__C (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__C (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A1 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__I1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A2 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__I (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__I (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__I (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__I (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__C (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__C (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__C (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__C (.I(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__I (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__I (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__C (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__C (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A4 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A4 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__C (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A3 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__I1 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A2 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A2 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__I (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__I (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__I (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__B (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__I (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__I (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A1 (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__I (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__C (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__C (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__C (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__C (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__C (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__C (.I(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__C (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__I (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__I (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__B2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__C (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__C (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__C (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__C (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__B (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__C (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__C1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__B (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__B (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__I (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__B (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__B (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__B (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__B (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A2 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__B2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__B2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__B (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__C (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__C (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__C (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__C (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__B (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__B (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__B (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__B (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A2 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A1 (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__I (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A2 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A2 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A4 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A3 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__B2 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A3 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A1 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A3 (.I(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A2 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__B2 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__B1 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__I (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A3 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__A1 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A4 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A1 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A4 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A3 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__I (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A1 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__B2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__I (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__I (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A2 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__B1 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__B2 (.I(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__B2 (.I(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__B1 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__B2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__I (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__B1 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__B2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A3 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A1 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A4 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A3 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A4 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__B2 (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__B (.I(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A2 (.I(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A2 (.I(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__I (.I(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__B (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__I (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A3 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__B1 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__B2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A3 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A2 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__B2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__B (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__B1 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__B2 (.I(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__C (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__C (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__C (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__C (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__S (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__I (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__I (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__I (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__B1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A2 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__I (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__I (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__I (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__B (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__B1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__I (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__I (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__I (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A2 (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A2 (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A2 (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__I (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__I (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__I (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__I (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__B1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__B1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__B1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__B1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__C (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__C (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__C (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__C (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A2 (.I(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__B1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__B1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__B1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__B1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__I (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__I (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__I (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__I (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__B (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__I (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__I (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__I (.I(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__I (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__I (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B1 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B1 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__B1 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__B1 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A2 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A2 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A2 (.I(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__B1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__B1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__B1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__I (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__I (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__I (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__I (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__B (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__B (.I(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__S (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__I (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__I (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__I (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A2 (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A2 (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__S (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__S (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A1 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A2 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A4 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__I (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__I (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__B1 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A3 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__I (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__B1 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__B1 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A2 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__B1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__B1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__I (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__I (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__I (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__I (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__I (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A2 (.I(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A1 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A2 (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A1 (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__I (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__B1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__B1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__I (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__I (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__B (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__B2 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__B2 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__I (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__I (.I(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__B (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__B (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__B (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__B (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__B (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__B (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__B (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A2 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A2 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A2 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A2 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__B (.I(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__B (.I(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__B (.I(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__B (.I(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__B1 (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__B1 (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__B1 (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A2 (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A2 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A2 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A2 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A2 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__I (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__B1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__B1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__B1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__B1 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__A1 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__B1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__I (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__I (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A2 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A1 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A2 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__B1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__B1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__B1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__B1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__B1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__B1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__B1 (.I(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A2 (.I(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A2 (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A2 (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__I (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A2 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A2 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A2 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__B1 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__B1 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__B1 (.I(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__B1 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__B1 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__B1 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__B1 (.I(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A2 (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A2 (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__I (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A2 (.I(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A2 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A2 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A2 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A2 (.I(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A2 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__B1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__B1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__B1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__B1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A2 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__B1 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__I (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__B1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__B1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__B1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__B1 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B1 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B1 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__B1 (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__B1 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__I (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__I (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A2 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A2 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__I (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__I (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A3 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__I (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__I (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A3 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A2 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A2 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__I (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A2 (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__B1 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__B1 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__B1 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clock_I (.I(clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(\cycles_per_ms[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__I (.I(\cycles_per_ms[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(\cycles_per_ms[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__I (.I(\cycles_per_ms[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__B2 (.I(\cycles_per_ms[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A1 (.I(\cycles_per_ms[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A1 (.I(\cycles_per_ms[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A4 (.I(\cycles_per_ms[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__I (.I(\cycles_per_ms[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(\delay_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A1 (.I(\delay_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A4 (.I(\delay_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(\delay_cycles[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(\delay_cycles[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(\delay_cycles[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__I (.I(\delay_cycles[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__B2 (.I(edge_interrupts));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(edge_interrupts));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__A1 (.I(edge_interrupts));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__I0 (.I(\exec.memory_input[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(\exec.memory_input[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I0 (.I(\exec.memory_input[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(\exec.memory_input[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I0 (.I(\exec.memory_input[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(\exec.memory_input[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__I0 (.I(\exec.memory_input[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(\exec.memory_input[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__I0 (.I(\exec.memory_input[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A1 (.I(\exec.memory_input[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(\exec.out_of_order_exec ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(\exec.out_of_order_exec ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(\exec.out_of_order_exec ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(i_la_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(i_la_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(i_la_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(i_la_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(i_la_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(i_la_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(i_la_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(i_la_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(i_la_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(i_la_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(i_la_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(i_la_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(i_la_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(i_la_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(i_la_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(i_la_wb_disable));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(i_la_write));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(i_wb_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(i_wb_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(i_wb_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(i_wb_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(i_wb_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(i_wb_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(i_wb_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(i_wb_addr[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(i_wb_addr[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(i_wb_addr[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(i_wb_addr[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(i_wb_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(i_wb_addr[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(i_wb_addr[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(i_wb_addr[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(i_wb_addr[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(i_wb_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(i_wb_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(i_wb_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(i_wb_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(i_wb_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(i_wb_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(i_wb_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(i_wb_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(i_wb_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(i_wb_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(i_wb_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(i_wb_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(i_wb_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(i_wb_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(i_wb_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(i_wb_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(i_wb_data[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(i_wb_data[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(i_wb_data[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(i_wb_data[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(i_wb_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(i_wb_data[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(i_wb_data[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(i_wb_data[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(i_wb_data[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(i_wb_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(i_wb_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(i_wb_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(i_wb_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(i_wb_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(i_wb_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(i_wb_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(i_wb_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(i_wb_stb));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(i_wb_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__B2 (.I(\intr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__B (.I(\intr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__A2 (.I(\intr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__B2 (.I(\intr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__B (.I(\intr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__B1 (.I(\intr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A2 (.I(\mem.dff_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__I0 (.I(\mem.dff_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(\mem.dff_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I0 (.I(\mem.dff_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(\mem.io_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(\mem.io_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__I0 (.I(\mem.io_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(\mem.io_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(\mem.io_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(\mem.io_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A1 (.I(\mem.mem_dff.code_mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I (.I(\mem.mem_dff.code_mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A1 (.I(\mem.mem_dff.code_mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__I (.I(\mem.mem_dff.code_mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(\mem.mem_dff.code_mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I (.I(\mem.mem_dff.code_mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(\mem.mem_dff.code_mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__I (.I(\mem.mem_dff.code_mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__B2 (.I(\mem.mem_dff.code_mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__I (.I(\mem.mem_dff.code_mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__B2 (.I(\mem.mem_dff.code_mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__I (.I(\mem.mem_dff.code_mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(\mem.mem_dff.code_mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__I (.I(\mem.mem_dff.code_mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__B2 (.I(\mem.mem_dff.code_mem[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__I (.I(\mem.mem_dff.code_mem[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__B2 (.I(\mem.mem_dff.code_mem[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__I (.I(\mem.mem_dff.code_mem[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__B2 (.I(\mem.mem_dff.code_mem[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__I (.I(\mem.mem_dff.code_mem[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__B2 (.I(\mem.mem_dff.code_mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(\mem.mem_dff.code_mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(\mem.mem_dff.code_mem[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__I (.I(\mem.mem_dff.code_mem[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__B2 (.I(\mem.mem_dff.code_mem[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__I (.I(\mem.mem_dff.code_mem[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__B2 (.I(\mem.mem_dff.code_mem[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__I (.I(\mem.mem_dff.code_mem[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(\mem.mem_dff.code_mem[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__I (.I(\mem.mem_dff.code_mem[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__B2 (.I(\mem.mem_dff.code_mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(\mem.mem_dff.code_mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__B2 (.I(\mem.mem_dff.code_mem[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(\mem.mem_dff.code_mem[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__B2 (.I(\mem.mem_dff.code_mem[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__I (.I(\mem.mem_dff.code_mem[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__B2 (.I(\mem.mem_dff.code_mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__I (.I(\mem.mem_dff.code_mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__B2 (.I(\mem.mem_dff.code_mem[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I (.I(\mem.mem_dff.code_mem[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__C1 (.I(\mem.mem_dff.code_mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__I (.I(\mem.mem_dff.code_mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(\mem.mem_dff.code_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I (.I(\mem.mem_dff.code_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(\mem.mem_dff.code_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__I (.I(\mem.mem_dff.code_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A1 (.I(\mem.mem_dff.code_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__I (.I(\mem.mem_dff.code_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(\mem.mem_dff.code_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__I (.I(\mem.mem_dff.code_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(\mem.mem_dff.code_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__I (.I(\mem.mem_dff.code_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(\mem.mem_dff.code_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I (.I(\mem.mem_dff.code_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(\mem.mem_dff.code_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__I (.I(\mem.mem_dff.code_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__B2 (.I(\mem.mem_dff.code_mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__I (.I(\mem.mem_dff.code_mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__B2 (.I(\mem.mem_dff.code_mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__I (.I(\mem.mem_dff.code_mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__B2 (.I(\mem.mem_dff.code_mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__I (.I(\mem.mem_dff.code_mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__C1 (.I(\mem.mem_dff.code_mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__I (.I(\mem.mem_dff.code_mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__C1 (.I(\mem.mem_dff.code_mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I (.I(\mem.mem_dff.code_mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__C1 (.I(\mem.mem_dff.code_mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__I (.I(\mem.mem_dff.code_mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__B2 (.I(\mem.mem_dff.code_mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(\mem.mem_dff.code_mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__B2 (.I(\mem.mem_dff.code_mem[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(\mem.mem_dff.code_mem[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__B2 (.I(\mem.mem_dff.code_mem[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(\mem.mem_dff.code_mem[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__B2 (.I(\mem.mem_dff.code_mem[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(\mem.mem_dff.code_mem[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__B2 (.I(\mem.mem_dff.code_mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(\mem.mem_dff.code_mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(\mem.mem_dff.code_mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(\mem.mem_dff.code_mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__B2 (.I(\mem.mem_dff.code_mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(\mem.mem_dff.code_mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(\mem.mem_dff.code_mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__I (.I(\mem.mem_dff.code_mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A1 (.I(\mem.mem_dff.code_mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(\mem.mem_dff.code_mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A1 (.I(\mem.mem_dff.code_mem[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__I (.I(\mem.mem_dff.code_mem[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(\mem.mem_dff.code_mem[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__I (.I(\mem.mem_dff.code_mem[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(\mem.mem_dff.code_mem[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__I (.I(\mem.mem_dff.code_mem[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(\mem.mem_dff.code_mem[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__I (.I(\mem.mem_dff.code_mem[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A1 (.I(\mem.mem_dff.code_mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__I (.I(\mem.mem_dff.code_mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A1 (.I(\mem.mem_dff.code_mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__I (.I(\mem.mem_dff.code_mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__A1 (.I(\mem.mem_dff.code_mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__I (.I(\mem.mem_dff.code_mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(\mem.mem_dff.code_mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__I (.I(\mem.mem_dff.code_mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A1 (.I(\mem.mem_dff.code_mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__I (.I(\mem.mem_dff.code_mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(\mem.mem_dff.code_mem[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__I (.I(\mem.mem_dff.code_mem[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__C1 (.I(\mem.mem_dff.code_mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(\mem.mem_dff.code_mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__C1 (.I(\mem.mem_dff.code_mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(\mem.mem_dff.code_mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__C1 (.I(\mem.mem_dff.code_mem[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__I (.I(\mem.mem_dff.code_mem[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__C1 (.I(\mem.mem_dff.code_mem[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__I (.I(\mem.mem_dff.code_mem[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__B2 (.I(\mem.mem_dff.code_mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(\mem.mem_dff.code_mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__B2 (.I(\mem.mem_dff.code_mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(\mem.mem_dff.code_mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__B2 (.I(\mem.mem_dff.code_mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__I (.I(\mem.mem_dff.code_mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__B2 (.I(\mem.mem_dff.code_mem[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I (.I(\mem.mem_dff.code_mem[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__B2 (.I(\mem.mem_dff.code_mem[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(\mem.mem_dff.code_mem[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__B2 (.I(\mem.mem_dff.code_mem[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__I (.I(\mem.mem_dff.code_mem[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__B2 (.I(\mem.mem_dff.code_mem[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__I (.I(\mem.mem_dff.code_mem[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(\mem.mem_dff.code_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(\mem.mem_dff.code_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(\mem.mem_dff.code_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__I (.I(\mem.mem_dff.code_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(\mem.mem_dff.code_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__I (.I(\mem.mem_dff.code_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(\mem.mem_dff.code_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__I (.I(\mem.mem_dff.code_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A1 (.I(\mem.mem_dff.code_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I (.I(\mem.mem_dff.code_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(\mem.mem_dff.code_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I (.I(\mem.mem_dff.code_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__C1 (.I(\mem.mem_dff.code_mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__I (.I(\mem.mem_dff.code_mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__C1 (.I(\mem.mem_dff.code_mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__I (.I(\mem.mem_dff.code_mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__B2 (.I(\mem.mem_dff.code_mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__I (.I(\mem.mem_dff.code_mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__B2 (.I(\mem.mem_dff.code_mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__I (.I(\mem.mem_dff.code_mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__C1 (.I(\mem.mem_dff.code_mem[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I (.I(\mem.mem_dff.code_mem[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__B2 (.I(\mem.mem_dff.code_mem[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__I (.I(\mem.mem_dff.code_mem[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__B2 (.I(\mem.mem_dff.code_mem[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__I (.I(\mem.mem_dff.code_mem[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__B2 (.I(\mem.mem_dff.code_mem[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__I (.I(\mem.mem_dff.code_mem[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A1 (.I(\mem.mem_dff.code_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__I (.I(\mem.mem_dff.code_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(\mem.mem_dff.code_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__I (.I(\mem.mem_dff.code_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A1 (.I(\mem.mem_dff.code_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__I (.I(\mem.mem_dff.code_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(\mem.mem_dff.code_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__I (.I(\mem.mem_dff.code_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(\mem.mem_dff.code_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__I (.I(\mem.mem_dff.code_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(\mem.mem_dff.code_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I (.I(\mem.mem_dff.code_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A1 (.I(\mem.mem_dff.code_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__I (.I(\mem.mem_dff.code_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(\mem.mem_dff.code_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I (.I(\mem.mem_dff.code_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(\mem.mem_dff.code_mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__I (.I(\mem.mem_dff.code_mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(\mem.mem_dff.code_mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__I (.I(\mem.mem_dff.code_mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(\mem.mem_dff.code_mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__I (.I(\mem.mem_dff.code_mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(\mem.mem_dff.code_mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__I (.I(\mem.mem_dff.code_mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(\mem.mem_dff.data_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__I (.I(\mem.mem_dff.data_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(\mem.mem_dff.data_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__I (.I(\mem.mem_dff.data_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A1 (.I(\mem.mem_dff.data_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__I (.I(\mem.mem_dff.data_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(\mem.mem_dff.data_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__I (.I(\mem.mem_dff.data_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A1 (.I(\mem.mem_dff.data_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__I (.I(\mem.mem_dff.data_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__B2 (.I(\mem.mem_dff.data_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(\mem.mem_dff.data_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__B2 (.I(\mem.mem_dff.data_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(\mem.mem_dff.data_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__B2 (.I(\mem.mem_dff.data_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__I (.I(\mem.mem_dff.data_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__B2 (.I(\mem.mem_dff.data_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__I (.I(\mem.mem_dff.data_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__B2 (.I(\mem.mem_dff.data_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(\mem.mem_dff.data_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__B2 (.I(\mem.mem_dff.data_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__I (.I(\mem.mem_dff.data_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__B2 (.I(\mem.mem_dff.data_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__I (.I(\mem.mem_dff.data_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__B2 (.I(\mem.mem_dff.data_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I (.I(\mem.mem_dff.data_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__C1 (.I(\mem.mem_dff.data_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A1 (.I(\mem.mem_dff.data_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__C1 (.I(\mem.mem_dff.data_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(\mem.mem_dff.data_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__C1 (.I(\mem.mem_dff.data_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A1 (.I(\mem.mem_dff.data_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__C1 (.I(\mem.mem_dff.data_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A1 (.I(\mem.mem_dff.data_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__I (.I(\mem.sram_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__I (.I(\mem.sram_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(rambus_wb_ack_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__CLK (.I(clknet_leaf_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(rambus_wb_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(rambus_wb_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(rambus_wb_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(rambus_wb_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(rambus_wb_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(rambus_wb_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(rambus_wb_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(rambus_wb_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(rambus_wb_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(rambus_wb_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(rambus_wb_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(rambus_wb_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(rambus_wb_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(rambus_wb_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(rambus_wb_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(rambus_wb_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(rambus_wb_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(rambus_wb_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(rambus_wb_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(rambus_wb_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(rambus_wb_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(rambus_wb_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(rambus_wb_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(rambus_wb_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(rambus_wb_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(rambus_wb_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(rambus_wb_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(rambus_wb_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(rambus_wb_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(rambus_wb_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(rambus_wb_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(rambus_wb_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(reset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(single_step));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A1 (.I(single_step));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__I (.I(single_step));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__B (.I(single_step));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__B2 (.I(\stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__I2 (.I(\stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__I1 (.I(\stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__B2 (.I(\stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I0 (.I(\stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__I1 (.I(\stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__B2 (.I(\stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__I2 (.I(\stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__I1 (.I(\stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__B2 (.I(\stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I0 (.I(\stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__A2 (.I(\stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__B2 (.I(\stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I2 (.I(\stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__A2 (.I(\stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__B2 (.I(\stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I2 (.I(\stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__A2 (.I(\stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__B2 (.I(\stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I2 (.I(\stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A2 (.I(\stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__B2 (.I(\stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I2 (.I(\stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A2 (.I(\stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__B2 (.I(\stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A2 (.I(\stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__I3 (.I(\stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__B2 (.I(\stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__I0 (.I(\stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__I3 (.I(\stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__B2 (.I(\stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__I0 (.I(\stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__I3 (.I(\stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__B2 (.I(\stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__I0 (.I(\stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__I3 (.I(\stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__B2 (.I(\stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__I0 (.I(\stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__I3 (.I(\stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__B2 (.I(\stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__I0 (.I(\stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__I3 (.I(\stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A1 (.I(\stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I0 (.I(\stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__B2 (.I(\stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(\stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__I0 (.I(\stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__B2 (.I(\stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(\stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__I1 (.I(\stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__I0 (.I(\stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__B2 (.I(\stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I1 (.I(\stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A2 (.I(\stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(\stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__I1 (.I(\stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__A2 (.I(\stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(\stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__I0 (.I(\stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__I1 (.I(\stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__B2 (.I(\stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I0 (.I(\stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__I1 (.I(\stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__B2 (.I(\stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__I0 (.I(\stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__I1 (.I(\stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__B2 (.I(\stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__I0 (.I(\stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__I1 (.I(\stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B2 (.I(\stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I0 (.I(\stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__A2 (.I(\stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__B2 (.I(\stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__I0 (.I(\stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A2 (.I(\stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(\stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__I1 (.I(\stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__I2 (.I(\stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__B2 (.I(\stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I1 (.I(\stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__I2 (.I(\stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__B2 (.I(\stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__I1 (.I(\stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__I2 (.I(\stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__B2 (.I(\stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I1 (.I(\stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__I2 (.I(\stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__B2 (.I(\stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__I1 (.I(\stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__I0 (.I(\stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__B2 (.I(\stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__I1 (.I(\stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__I0 (.I(\stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__B2 (.I(\stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I1 (.I(\stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__B1 (.I(\stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(\stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__I1 (.I(\stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__B1 (.I(\stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__B2 (.I(\stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__A2 (.I(\stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__I3 (.I(\stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__B2 (.I(\stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I0 (.I(\stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__I3 (.I(\stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__B2 (.I(\stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__I0 (.I(\stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__I3 (.I(\stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__B2 (.I(\stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__I0 (.I(\stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__I3 (.I(\stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__B2 (.I(\stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__I0 (.I(\stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__A1 (.I(\stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__B2 (.I(\stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__I0 (.I(\stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__A1 (.I(\stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(\stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I0 (.I(\stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__A1 (.I(\stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__B2 (.I(\stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__I0 (.I(\stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__A1 (.I(\stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__I (.I(\stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__I0 (.I(\stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__I (.I(\stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I1 (.I(\stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__I0 (.I(\stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__I (.I(\stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__I1 (.I(\stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__I0 (.I(\stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__I (.I(\stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__I1 (.I(\stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__I0 (.I(\stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__I (.I(\stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__I1 (.I(\stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05443__A1 (.I(\stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__B2 (.I(\stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__I1 (.I(\stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__A1 (.I(\stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__B2 (.I(\stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I1 (.I(\stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__B2 (.I(\stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__B2 (.I(\stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__I1 (.I(\stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__B2 (.I(\stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__B2 (.I(\stack[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I2 (.I(\stack[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__I1 (.I(\stack[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B2 (.I(\stack[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I2 (.I(\stack[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A2 (.I(\stack[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B2 (.I(\stack[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I2 (.I(\stack[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__A2 (.I(\stack[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__B2 (.I(\stack[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I3 (.I(\stack[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__I2 (.I(\stack[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B2 (.I(\stack[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I3 (.I(\stack[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__B1 (.I(\stack[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(\stack[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__I1 (.I(\stack[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__B1 (.I(\stack[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__B2 (.I(\stack[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I0 (.I(\stack[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__I3 (.I(\stack[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__B2 (.I(\stack[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I0 (.I(\stack[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__I3 (.I(\stack[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__B2 (.I(\stack[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I0 (.I(\stack[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__I3 (.I(\stack[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__B2 (.I(\stack[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__I0 (.I(\stack[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__I3 (.I(\stack[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__B2 (.I(\stack[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__I0 (.I(\stack[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__B2 (.I(\stack[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__B2 (.I(\stack[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I0 (.I(\stack[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__B2 (.I(\stack[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(\stack[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I0 (.I(\stack[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__B2 (.I(\stack[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__B2 (.I(\stack[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__I0 (.I(\stack[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__A1 (.I(\stack[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__B2 (.I(\stack[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I1 (.I(\stack[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__I0 (.I(\stack[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__B2 (.I(\stack[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I1 (.I(\stack[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__I0 (.I(\stack[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__B2 (.I(\stack[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I1 (.I(\stack[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__I0 (.I(\stack[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__B2 (.I(\stack[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__I1 (.I(\stack[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__I0 (.I(\stack[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__B2 (.I(\stack[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__I1 (.I(\stack[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__A2 (.I(\stack[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__B2 (.I(\stack[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I1 (.I(\stack[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__A2 (.I(\stack[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__B2 (.I(\stack[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I1 (.I(\stack[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__A2 (.I(\stack[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__B2 (.I(\stack[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__I1 (.I(\stack[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__B2 (.I(\stack[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(\stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__I3 (.I(\stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__I2 (.I(\stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__B2 (.I(\stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I1 (.I(\stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__I2 (.I(\stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__B2 (.I(\stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__I3 (.I(\stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__I2 (.I(\stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__B2 (.I(\stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__I1 (.I(\stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__B1 (.I(\stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__B2 (.I(\stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I3 (.I(\stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__B1 (.I(\stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__B2 (.I(\stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I3 (.I(\stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__B1 (.I(\stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__B2 (.I(\stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I3 (.I(\stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__B1 (.I(\stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__B2 (.I(\stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I3 (.I(\stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__B1 (.I(\stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A1 (.I(\stack[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I0 (.I(\stack[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__I1 (.I(\stack[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__B2 (.I(\stack[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I0 (.I(\stack[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__I1 (.I(\stack[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__B2 (.I(\stack[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__I0 (.I(\stack[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__I1 (.I(\stack[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__B2 (.I(\stack[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I0 (.I(\stack[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__A2 (.I(\stack[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__B2 (.I(\stack[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(\stack[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__A2 (.I(\stack[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__B2 (.I(\stack[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I0 (.I(\stack[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__I1 (.I(\stack[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__B2 (.I(\stack[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__I0 (.I(\stack[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__I1 (.I(\stack[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__B2 (.I(\stack[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I0 (.I(\stack[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__A2 (.I(\stack[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(\stack[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I1 (.I(\stack[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__I2 (.I(\stack[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__B2 (.I(\stack[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I1 (.I(\stack[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__I2 (.I(\stack[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__B2 (.I(\stack[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__I1 (.I(\stack[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__I2 (.I(\stack[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__B2 (.I(\stack[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I1 (.I(\stack[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__B1 (.I(\stack[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__B2 (.I(\stack[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A2 (.I(\stack[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__B1 (.I(\stack[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__B2 (.I(\stack[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I1 (.I(\stack[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__I2 (.I(\stack[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__B2 (.I(\stack[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__I1 (.I(\stack[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__I2 (.I(\stack[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A1 (.I(\stack[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I1 (.I(\stack[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__B1 (.I(\stack[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__B2 (.I(\stack[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__I0 (.I(\stack[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__I3 (.I(\stack[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__B2 (.I(\stack[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I0 (.I(\stack[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__I3 (.I(\stack[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__B2 (.I(\stack[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__I0 (.I(\stack[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__I3 (.I(\stack[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__B2 (.I(\stack[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I0 (.I(\stack[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A3 (.I(\stack[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__B2 (.I(\stack[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__A2 (.I(\stack[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__A1 (.I(\stack[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A1 (.I(\stack[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I0 (.I(\stack[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__I3 (.I(\stack[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__B2 (.I(\stack[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I0 (.I(\stack[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__A1 (.I(\stack[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(\stack[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I1 (.I(\stack[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__I0 (.I(\stack[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(\stack[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I1 (.I(\stack[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__A1 (.I(\stack[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(\stack[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A2 (.I(\stack[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__B2 (.I(\stack[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__B2 (.I(\stack[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I1 (.I(\stack[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__I0 (.I(\stack[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(\stack[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I1 (.I(\stack[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__B2 (.I(\stack[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__B2 (.I(\stack[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__I0 (.I(\stack[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__I1 (.I(\stack[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__B2 (.I(\stack[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__I0 (.I(\stack[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__I1 (.I(\stack[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__B2 (.I(\stack[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__I0 (.I(\stack[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__I1 (.I(\stack[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__B2 (.I(\stack[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I0 (.I(\stack[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__I1 (.I(\stack[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__B2 (.I(\stack[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I0 (.I(\stack[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__I1 (.I(\stack[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__B2 (.I(\stack[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__I0 (.I(\stack[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__A2 (.I(\stack[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__B2 (.I(\stack[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I0 (.I(\stack[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__A2 (.I(\stack[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(\stack[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__I0 (.I(\stack[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__A2 (.I(\stack[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(\stack[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__I1 (.I(\stack[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__I2 (.I(\stack[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__B2 (.I(\stack[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__I1 (.I(\stack[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__I2 (.I(\stack[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__B2 (.I(\stack[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__I1 (.I(\stack[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__I2 (.I(\stack[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__B2 (.I(\stack[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I1 (.I(\stack[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__I2 (.I(\stack[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__B2 (.I(\stack[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I1 (.I(\stack[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__I2 (.I(\stack[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__B2 (.I(\stack[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__I1 (.I(\stack[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__B1 (.I(\stack[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__B2 (.I(\stack[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I1 (.I(\stack[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__B1 (.I(\stack[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(\stack[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__I1 (.I(\stack[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__B1 (.I(\stack[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__B2 (.I(\stack[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__I0 (.I(\stack[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__I3 (.I(\stack[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B2 (.I(\stack[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__I0 (.I(\stack[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__I3 (.I(\stack[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__B2 (.I(\stack[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__A2 (.I(\stack[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__I3 (.I(\stack[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__B2 (.I(\stack[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I0 (.I(\stack[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__I3 (.I(\stack[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__B2 (.I(\stack[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__I0 (.I(\stack[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__I3 (.I(\stack[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__B2 (.I(\stack[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I0 (.I(\stack[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__A1 (.I(\stack[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(\stack[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__I0 (.I(\stack[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__B2 (.I(\stack[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(\stack[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__I0 (.I(\stack[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__B2 (.I(\stack[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(\stack[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__A2 (.I(\stack[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__I0 (.I(\stack[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(\stack[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I1 (.I(\stack[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__B2 (.I(\stack[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__B2 (.I(\stack[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__I1 (.I(\stack[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__A2 (.I(\stack[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(\stack[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__I1 (.I(\stack[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__A2 (.I(\stack[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(\stack[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__I0 (.I(\stack[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__I1 (.I(\stack[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__B2 (.I(\stack[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I0 (.I(\stack[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__I1 (.I(\stack[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__B2 (.I(\stack[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__I0 (.I(\stack[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__I1 (.I(\stack[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__B2 (.I(\stack[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I0 (.I(\stack[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__I1 (.I(\stack[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__B2 (.I(\stack[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__I0 (.I(\stack[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__A2 (.I(\stack[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__B2 (.I(\stack[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I0 (.I(\stack[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__A2 (.I(\stack[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B2 (.I(\stack[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I0 (.I(\stack[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__A2 (.I(\stack[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__B2 (.I(\stack[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__I0 (.I(\stack[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__A2 (.I(\stack[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B2 (.I(\stack[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I1 (.I(\stack[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__I2 (.I(\stack[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__B2 (.I(\stack[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__I1 (.I(\stack[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__I2 (.I(\stack[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__B2 (.I(\stack[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I1 (.I(\stack[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__I2 (.I(\stack[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__B2 (.I(\stack[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__I1 (.I(\stack[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__B1 (.I(\stack[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B2 (.I(\stack[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I1 (.I(\stack[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__B1 (.I(\stack[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__B2 (.I(\stack[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I1 (.I(\stack[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__B1 (.I(\stack[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__B2 (.I(\stack[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__I1 (.I(\stack[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__B1 (.I(\stack[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(\stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I0 (.I(\stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__I3 (.I(\stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(\stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__I0 (.I(\stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__I3 (.I(\stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A1 (.I(\stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I0 (.I(\stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__B2 (.I(\stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(\stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I0 (.I(\stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__B2 (.I(\stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A1 (.I(\stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I0 (.I(\stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__B2 (.I(\stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__B2 (.I(\stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I0 (.I(\stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__B2 (.I(\stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__B2 (.I(\stack[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I0 (.I(\stack[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__I3 (.I(\stack[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__B2 (.I(\stack[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__I0 (.I(\stack[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A1 (.I(\stack[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__B2 (.I(\stack[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__I0 (.I(\stack[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__A1 (.I(\stack[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(\stack[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__I0 (.I(\stack[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A1 (.I(\stack[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__I (.I(\stack[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__I0 (.I(\stack[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__I (.I(\stack[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I1 (.I(\stack[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__I0 (.I(\stack[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__I (.I(\stack[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__I0 (.I(\stack[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__I (.I(\stack[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I1 (.I(\stack[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__I0 (.I(\stack[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__I (.I(\stack[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__I1 (.I(\stack[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__B2 (.I(\stack[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(\stack[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__I1 (.I(\stack[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__B2 (.I(\stack[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(\stack[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__I1 (.I(\stack[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__B2 (.I(\stack[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(\stack[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__I1 (.I(\stack[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__B2 (.I(\stack[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A1 (.I(\stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I1 (.I(\stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__I0 (.I(\stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A1 (.I(\stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__I1 (.I(\stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__A2 (.I(\stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(\stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I1 (.I(\stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__A2 (.I(\stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__B2 (.I(\stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I1 (.I(\stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__A2 (.I(\stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__B2 (.I(\stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I1 (.I(\stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A2 (.I(\stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__B2 (.I(\stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I1 (.I(\stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__A2 (.I(\stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B2 (.I(\stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A2 (.I(\stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__I1 (.I(\stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__B2 (.I(\stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A2 (.I(\stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__A2 (.I(\stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__B2 (.I(\stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I0 (.I(\stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__A2 (.I(\stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__B2 (.I(\stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__I0 (.I(\stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__I1 (.I(\stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(\stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__I1 (.I(\stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__I2 (.I(\stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__B2 (.I(\stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__I1 (.I(\stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__I2 (.I(\stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B2 (.I(\stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A2 (.I(\stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__I2 (.I(\stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B2 (.I(\stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__I1 (.I(\stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__I0 (.I(\stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__B2 (.I(\stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A2 (.I(\stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__B1 (.I(\stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B2 (.I(\stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I1 (.I(\stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__B1 (.I(\stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B2 (.I(\stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__I1 (.I(\stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__I2 (.I(\stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(\stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__I0 (.I(\stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__I3 (.I(\stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B2 (.I(\stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A2 (.I(\stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A1 (.I(\stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A1 (.I(\stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__I0 (.I(\stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__A1 (.I(\stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(\stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I0 (.I(\stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__I3 (.I(\stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(\stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__I1 (.I(\stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__I0 (.I(\stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A1 (.I(\stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I1 (.I(\stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__I0 (.I(\stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(\stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__A2 (.I(\stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__I0 (.I(\stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A1 (.I(\stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__I1 (.I(\stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__A1 (.I(\stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(\stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A2 (.I(\stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__B2 (.I(\stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B2 (.I(\stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__I1 (.I(\stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__I0 (.I(\stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__B2 (.I(\stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__I1 (.I(\stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__A1 (.I(\stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__B2 (.I(\stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I1 (.I(\stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__I0 (.I(\stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__B2 (.I(\stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__I0 (.I(\stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__I1 (.I(\stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__B2 (.I(\stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__I0 (.I(\stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__I1 (.I(\stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__B2 (.I(\stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__I1 (.I(\stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__I2 (.I(\stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__B2 (.I(\stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I1 (.I(\stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__I2 (.I(\stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__B2 (.I(\stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__I1 (.I(\stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__I2 (.I(\stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__B2 (.I(\stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__I1 (.I(\stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__I2 (.I(\stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B2 (.I(\stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__I1 (.I(\stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__I2 (.I(\stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__B2 (.I(\stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__I1 (.I(\stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__I2 (.I(\stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__B2 (.I(\stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__I1 (.I(\stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__B1 (.I(\stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(\stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__I1 (.I(\stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__B1 (.I(\stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__S (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__B (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A4 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A3 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A4 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A3 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A4 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A4 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A3 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I0 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I0 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__I0 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__I0 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A3 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__B2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__B2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__B2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__B2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__B2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__B2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__B2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__B2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__B2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__B2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__B2 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__B2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__B2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__B2 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__B2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A2 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__B2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__B2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__B2 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__B2 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__B2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__B2 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__B2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__B2 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__B2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__B2 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__B2 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__B2 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__B2 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__C2 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__B2 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__B2 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__B2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__B2 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__B2 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__B2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B2 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__B2 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__B2 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__A2 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__A1 (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05646__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A4 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05641__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A3 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__A2 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05230__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05211__I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05231__I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05219__I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05218__I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A2 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05296__I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05223__I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__A1 (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output141_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A3 (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B2 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__B2 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__B2 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__B2 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__B2 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__B2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__B2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__B2 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__B2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__B2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__B2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A1 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__B2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__B2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout257_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__C1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A2 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A1 (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A1 (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A1 (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A1 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A1 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout255_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout254_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A2 (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05626__I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A1 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A2 (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__C (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A1 (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output194_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output195_I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A2 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A2 (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__C1 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A2 (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output229_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__B1 (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A2 (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout233_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout247_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout250_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout251_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output232_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A1 (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A1 (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output142_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__C1 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A1 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A1 (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A1 (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__CLK (.I(clknet_leaf_3_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__CLK (.I(clknet_leaf_5_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__CLK (.I(clknet_leaf_8_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__CLK (.I(clknet_leaf_9_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__CLK (.I(clknet_leaf_13_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__CLK (.I(clknet_leaf_14_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__CLK (.I(clknet_leaf_16_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__CLK (.I(clknet_leaf_17_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__CLK (.I(clknet_leaf_19_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__CLK (.I(clknet_leaf_25_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__CLK (.I(clknet_leaf_26_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__CLK (.I(clknet_leaf_29_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__CLK (.I(clknet_leaf_30_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__CLK (.I(clknet_leaf_31_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__CLK (.I(clknet_leaf_33_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__CLK (.I(clknet_leaf_34_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__CLK (.I(clknet_leaf_35_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__CLK (.I(clknet_leaf_36_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__CLK (.I(clknet_leaf_37_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__CLK (.I(clknet_leaf_38_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__CLK (.I(clknet_leaf_39_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__CLK (.I(clknet_leaf_40_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__CLK (.I(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__CLK (.I(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__CLK (.I(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__CLK (.I(clknet_leaf_41_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__CLK (.I(clknet_leaf_42_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__CLK (.I(clknet_leaf_43_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__CLK (.I(clknet_leaf_45_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__CLK (.I(clknet_leaf_45_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__CLK (.I(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__CLK (.I(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__CLK (.I(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__CLK (.I(clknet_leaf_48_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__CLK (.I(clknet_leaf_49_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__CLK (.I(clknet_leaf_50_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__CLK (.I(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__CLK (.I(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__CLK (.I(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__CLK (.I(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__CLK (.I(clknet_leaf_51_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__CLK (.I(clknet_leaf_53_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__CLK (.I(clknet_leaf_54_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__CLK (.I(clknet_leaf_55_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__CLK (.I(clknet_leaf_56_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__CLK (.I(clknet_leaf_57_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__CLK (.I(clknet_leaf_59_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__CLK (.I(clknet_leaf_60_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__CLK (.I(clknet_leaf_61_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__CLK (.I(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__CLK (.I(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__CLK (.I(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__CLK (.I(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__CLK (.I(clknet_leaf_62_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__CLK (.I(clknet_leaf_64_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__CLK (.I(clknet_leaf_67_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__CLK (.I(clknet_leaf_68_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__CLK (.I(clknet_leaf_69_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__CLK (.I(clknet_leaf_70_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__CLK (.I(clknet_leaf_72_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__CLK (.I(clknet_leaf_73_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__CLK (.I(clknet_leaf_75_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__CLK (.I(clknet_leaf_76_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__CLK (.I(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__CLK (.I(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__CLK (.I(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__CLK (.I(clknet_leaf_79_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__CLK (.I(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__CLK (.I(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__CLK (.I(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__CLK (.I(clknet_leaf_81_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__CLK (.I(clknet_leaf_82_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__CLK (.I(clknet_leaf_85_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__CLK (.I(clknet_leaf_86_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__CLK (.I(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__CLK (.I(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__CLK (.I(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__CLK (.I(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__CLK (.I(clknet_leaf_87_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__CLK (.I(clknet_leaf_89_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__CLK (.I(clknet_leaf_89_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__CLK (.I(clknet_leaf_89_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__CLK (.I(clknet_leaf_90_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__CLK (.I(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__CLK (.I(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__CLK (.I(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__CLK (.I(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__CLK (.I(clknet_leaf_92_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__CLK (.I(clknet_leaf_94_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__CLK (.I(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__CLK (.I(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__CLK (.I(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__CLK (.I(clknet_leaf_95_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__CLK (.I(clknet_leaf_96_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__CLK (.I(clknet_leaf_97_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__CLK (.I(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__CLK (.I(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__CLK (.I(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__CLK (.I(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__CLK (.I(clknet_leaf_99_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__CLK (.I(clknet_leaf_100_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__CLK (.I(clknet_leaf_101_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__CLK (.I(clknet_leaf_102_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__CLK (.I(clknet_leaf_103_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__CLK (.I(clknet_leaf_104_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__CLK (.I(clknet_leaf_105_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__CLK (.I(clknet_leaf_106_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__CLK (.I(clknet_leaf_107_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__CLK (.I(clknet_leaf_107_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__CLK (.I(clknet_leaf_107_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__CLK (.I(clknet_leaf_108_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__CLK (.I(clknet_leaf_110_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__CLK (.I(clknet_leaf_112_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__CLK (.I(clknet_leaf_113_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__CLK (.I(clknet_leaf_115_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__CLK (.I(clknet_leaf_116_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__CLK (.I(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__CLK (.I(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__CLK (.I(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__CLK (.I(clknet_leaf_117_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__CLK (.I(clknet_leaf_120_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__CLK (.I(clknet_leaf_122_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__CLK (.I(clknet_leaf_123_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__CLK (.I(clknet_leaf_125_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__CLK (.I(clknet_leaf_127_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__CLK (.I(clknet_leaf_128_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__CLK (.I(clknet_leaf_129_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__CLK (.I(clknet_leaf_135_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__CLK (.I(clknet_leaf_138_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__CLK (.I(clknet_leaf_139_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__CLK (.I(clknet_leaf_141_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__CLK (.I(clknet_leaf_142_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__CLK (.I(clknet_leaf_142_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__CLK (.I(clknet_leaf_142_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__CLK (.I(clknet_leaf_142_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__CLK (.I(clknet_leaf_143_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__CLK (.I(clknet_leaf_147_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__CLK (.I(clknet_leaf_148_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__CLK (.I(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__CLK (.I(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__CLK (.I(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__CLK (.I(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__CLK (.I(clknet_leaf_149_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__CLK (.I(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__CLK (.I(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__CLK (.I(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__CLK (.I(clknet_leaf_153_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__CLK (.I(clknet_leaf_158_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__CLK (.I(clknet_leaf_159_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__CLK (.I(clknet_leaf_160_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__CLK (.I(clknet_leaf_161_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__CLK (.I(clknet_leaf_162_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__CLK (.I(clknet_leaf_163_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__CLK (.I(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__CLK (.I(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__CLK (.I(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__CLK (.I(clknet_leaf_167_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__CLK (.I(clknet_leaf_168_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__CLK (.I(clknet_leaf_169_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__CLK (.I(clknet_leaf_170_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__CLK (.I(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__CLK (.I(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__CLK (.I(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__CLK (.I(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__CLK (.I(clknet_leaf_171_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__CLK (.I(clknet_leaf_173_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__CLK (.I(clknet_leaf_176_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__CLK (.I(clknet_leaf_176_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__CLK (.I(clknet_leaf_177_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__CLK (.I(clknet_leaf_177_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__CLK (.I(clknet_leaf_177_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__CLK (.I(clknet_leaf_178_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__CLK (.I(clknet_leaf_179_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__CLK (.I(clknet_leaf_180_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__CLK (.I(clknet_leaf_181_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__CLK (.I(clknet_leaf_183_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__CLK (.I(clknet_leaf_186_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__CLK (.I(clknet_leaf_187_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__CLK (.I(clknet_leaf_189_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__CLK (.I(clknet_leaf_190_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__CLK (.I(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__CLK (.I(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__CLK (.I(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__CLK (.I(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__CLK (.I(clknet_leaf_191_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__CLK (.I(clknet_leaf_192_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0_0_clock_I (.I(clknet_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_clock_I (.I(clknet_2_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_clock_I (.I(clknet_2_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_clock_I (.I(clknet_2_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_clock_I (.I(clknet_2_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_clock_I (.I(clknet_2_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_clock_I (.I(clknet_2_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_clock_I (.I(clknet_2_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_clock_I (.I(clknet_2_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_clock_I (.I(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_clock_I (.I(clknet_3_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_clock_I (.I(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_clock_I (.I(clknet_3_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_clock_I (.I(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_clock_I (.I(clknet_3_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_clock_I (.I(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_clock_I (.I(clknet_3_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_clock_I (.I(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_clock_I (.I(clknet_3_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_clock_I (.I(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_clock_I (.I(clknet_3_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_clock_I (.I(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_clock_I (.I(clknet_3_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_clock_I (.I(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_clock_I (.I(clknet_3_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__CLK (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_191_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__CLK (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clock_I (.I(clknet_4_0_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_193_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_192_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_190_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_189_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_188_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_187_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_186_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__CLK (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_173_clock_I (.I(clknet_4_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__CLK (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_clock_I (.I(clknet_4_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__CLK (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_171_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_170_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_169_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_168_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_167_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__CLK (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__CLK (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__CLK (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clock_I (.I(clknet_4_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_185_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_184_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_183_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_182_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_181_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_180_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_179_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_178_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_177_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_176_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_175_clock_I (.I(clknet_4_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_clock_I (.I(clknet_4_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clock_I (.I(clknet_4_6_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__CLK (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_clock_I (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__CLK (.I(clknet_4_7_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__CLK (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clock_I (.I(clknet_4_8_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__CLK (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__CLK (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clock_I (.I(clknet_4_9_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_4_0_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clock_I (.I(clknet_4_10_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_5_0_clock_I (.I(clknet_4_11_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_6_0_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__CLK (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__CLK (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clock_I (.I(clknet_4_12_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clock_I (.I(clknet_4_13_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__CLK (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clock_I (.I(clknet_4_14_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__CLK (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clock_I (.I(clknet_4_15_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__CLK (.I(clknet_opt_1_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__CLK (.I(clknet_opt_2_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__CLK (.I(clknet_opt_3_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_4_1_clock_I (.I(clknet_opt_4_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__I (.I(clknet_opt_4_1_clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__CLK (.I(clknet_opt_5_0_clock));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1577 ();
 assign o_wb_data[24] = net259;
 assign o_wb_data[25] = net260;
 assign o_wb_data[26] = net261;
 assign o_wb_data[27] = net262;
 assign o_wb_data[28] = net263;
 assign o_wb_data[29] = net264;
 assign o_wb_data[30] = net265;
 assign o_wb_data[31] = net266;
 assign rambus_wb_addr_o[0] = net267;
 assign rambus_wb_addr_o[1] = net268;
 assign rambus_wb_addr_o[9] = net269;
endmodule

