magic
tech gf180mcuC
magscale 1 5
timestamp 1670238422
<< obsm1 >>
rect 672 1538 279328 178457
<< metal2 >>
rect 8400 179600 8456 179900
rect 19488 179600 19544 179900
rect 30576 179600 30632 179900
rect 41664 179600 41720 179900
rect 52752 179600 52808 179900
rect 63840 179600 63896 179900
rect 74928 179600 74984 179900
rect 86016 179600 86072 179900
rect 97104 179600 97160 179900
rect 108192 179600 108248 179900
rect 119280 179600 119336 179900
rect 130368 179600 130424 179900
rect 141456 179600 141512 179900
rect 152544 179600 152600 179900
rect 163632 179600 163688 179900
rect 174720 179600 174776 179900
rect 185808 179600 185864 179900
rect 196896 179600 196952 179900
rect 207984 179600 208040 179900
rect 219072 179600 219128 179900
rect 230160 179600 230216 179900
rect 241248 179600 241304 179900
rect 252336 179600 252392 179900
rect 263424 179600 263480 179900
rect 274512 179600 274568 179900
rect 0 100 56 400
rect 11088 100 11144 400
rect 22176 100 22232 400
rect 33264 100 33320 400
rect 44352 100 44408 400
rect 55440 100 55496 400
rect 66528 100 66584 400
rect 77616 100 77672 400
rect 88704 100 88760 400
rect 99792 100 99848 400
rect 110880 100 110936 400
rect 121968 100 122024 400
rect 133056 100 133112 400
rect 144144 100 144200 400
rect 155232 100 155288 400
rect 166320 100 166376 400
rect 177408 100 177464 400
rect 188496 100 188552 400
rect 199584 100 199640 400
rect 210672 100 210728 400
rect 221760 100 221816 400
rect 232848 100 232904 400
rect 243936 100 243992 400
rect 255024 100 255080 400
rect 266112 100 266168 400
rect 277200 100 277256 400
<< obsm2 >>
rect 14 179930 279090 179970
rect 14 179570 8370 179930
rect 8486 179570 19458 179930
rect 19574 179570 30546 179930
rect 30662 179570 41634 179930
rect 41750 179570 52722 179930
rect 52838 179570 63810 179930
rect 63926 179570 74898 179930
rect 75014 179570 85986 179930
rect 86102 179570 97074 179930
rect 97190 179570 108162 179930
rect 108278 179570 119250 179930
rect 119366 179570 130338 179930
rect 130454 179570 141426 179930
rect 141542 179570 152514 179930
rect 152630 179570 163602 179930
rect 163718 179570 174690 179930
rect 174806 179570 185778 179930
rect 185894 179570 196866 179930
rect 196982 179570 207954 179930
rect 208070 179570 219042 179930
rect 219158 179570 230130 179930
rect 230246 179570 241218 179930
rect 241334 179570 252306 179930
rect 252422 179570 263394 179930
rect 263510 179570 274482 179930
rect 274598 179570 279090 179930
rect 14 430 279090 179570
rect 86 289 11058 430
rect 11174 289 22146 430
rect 22262 289 33234 430
rect 33350 289 44322 430
rect 44438 289 55410 430
rect 55526 289 66498 430
rect 66614 289 77586 430
rect 77702 289 88674 430
rect 88790 289 99762 430
rect 99878 289 110850 430
rect 110966 289 121938 430
rect 122054 289 133026 430
rect 133142 289 144114 430
rect 144230 289 155202 430
rect 155318 289 166290 430
rect 166406 289 177378 430
rect 177494 289 188466 430
rect 188582 289 199554 430
rect 199670 289 210642 430
rect 210758 289 221730 430
rect 221846 289 232818 430
rect 232934 289 243906 430
rect 244022 289 254994 430
rect 255110 289 266082 430
rect 266198 289 277170 430
rect 277286 289 279090 430
<< metal3 >>
rect 100 177408 400 177464
rect 279600 174384 279900 174440
rect 100 166320 400 166376
rect 279600 163296 279900 163352
rect 100 155232 400 155288
rect 279600 152208 279900 152264
rect 100 144144 400 144200
rect 279600 141120 279900 141176
rect 100 133056 400 133112
rect 279600 130032 279900 130088
rect 100 121968 400 122024
rect 279600 118944 279900 119000
rect 100 110880 400 110936
rect 279600 107856 279900 107912
rect 100 99792 400 99848
rect 279600 96768 279900 96824
rect 100 88704 400 88760
rect 279600 85680 279900 85736
rect 100 77616 400 77672
rect 279600 74592 279900 74648
rect 100 66528 400 66584
rect 279600 63504 279900 63560
rect 100 55440 400 55496
rect 279600 52416 279900 52472
rect 100 44352 400 44408
rect 279600 41328 279900 41384
rect 100 33264 400 33320
rect 279600 30240 279900 30296
rect 100 22176 400 22232
rect 279600 19152 279900 19208
rect 100 11088 400 11144
rect 279600 8064 279900 8120
<< obsm3 >>
rect 9 177494 279600 179690
rect 9 177378 70 177494
rect 430 177378 279600 177494
rect 9 174470 279600 177378
rect 9 174354 279570 174470
rect 9 166406 279600 174354
rect 9 166290 70 166406
rect 430 166290 279600 166406
rect 9 163382 279600 166290
rect 9 163266 279570 163382
rect 9 155318 279600 163266
rect 9 155202 70 155318
rect 430 155202 279600 155318
rect 9 152294 279600 155202
rect 9 152178 279570 152294
rect 9 144230 279600 152178
rect 9 144114 70 144230
rect 430 144114 279600 144230
rect 9 141206 279600 144114
rect 9 141090 279570 141206
rect 9 133142 279600 141090
rect 9 133026 70 133142
rect 430 133026 279600 133142
rect 9 130118 279600 133026
rect 9 130002 279570 130118
rect 9 122054 279600 130002
rect 9 121938 70 122054
rect 430 121938 279600 122054
rect 9 119030 279600 121938
rect 9 118914 279570 119030
rect 9 110966 279600 118914
rect 9 110850 70 110966
rect 430 110850 279600 110966
rect 9 107942 279600 110850
rect 9 107826 279570 107942
rect 9 99878 279600 107826
rect 9 99762 70 99878
rect 430 99762 279600 99878
rect 9 96854 279600 99762
rect 9 96738 279570 96854
rect 9 88790 279600 96738
rect 9 88674 70 88790
rect 430 88674 279600 88790
rect 9 85766 279600 88674
rect 9 85650 279570 85766
rect 9 77702 279600 85650
rect 9 77586 70 77702
rect 430 77586 279600 77702
rect 9 74678 279600 77586
rect 9 74562 279570 74678
rect 9 66614 279600 74562
rect 9 66498 70 66614
rect 430 66498 279600 66614
rect 9 63590 279600 66498
rect 9 63474 279570 63590
rect 9 55526 279600 63474
rect 9 55410 70 55526
rect 430 55410 279600 55526
rect 9 52502 279600 55410
rect 9 52386 279570 52502
rect 9 44438 279600 52386
rect 9 44322 70 44438
rect 430 44322 279600 44438
rect 9 41414 279600 44322
rect 9 41298 279570 41414
rect 9 33350 279600 41298
rect 9 33234 70 33350
rect 430 33234 279600 33350
rect 9 30326 279600 33234
rect 9 30210 279570 30326
rect 9 22262 279600 30210
rect 9 22146 70 22262
rect 430 22146 279600 22262
rect 9 19238 279600 22146
rect 9 19122 279570 19238
rect 9 11174 279600 19122
rect 9 11058 70 11174
rect 430 11058 279600 11174
rect 9 8150 279600 11058
rect 9 8034 279570 8150
rect 9 294 279600 8034
<< metal4 >>
rect 2224 1538 2384 178390
rect 9904 1538 10064 178390
rect 17584 1538 17744 178390
rect 25264 1538 25424 178390
rect 32944 1538 33104 178390
rect 40624 1538 40784 178390
rect 48304 1538 48464 178390
rect 55984 1538 56144 178390
rect 63664 1538 63824 178390
rect 71344 1538 71504 178390
rect 79024 1538 79184 178390
rect 86704 1538 86864 178390
rect 94384 1538 94544 178390
rect 102064 1538 102224 178390
rect 109744 1538 109904 178390
rect 117424 1538 117584 178390
rect 125104 1538 125264 178390
rect 132784 1538 132944 178390
rect 140464 1538 140624 178390
rect 148144 1538 148304 178390
rect 155824 1538 155984 178390
rect 163504 1538 163664 178390
rect 171184 1538 171344 178390
rect 178864 1538 179024 178390
rect 186544 1538 186704 178390
rect 194224 1538 194384 178390
rect 201904 1538 202064 178390
rect 209584 1538 209744 178390
rect 217264 1538 217424 178390
rect 224944 1538 225104 178390
rect 232624 1538 232784 178390
rect 240304 1538 240464 178390
rect 247984 1538 248144 178390
rect 255664 1538 255824 178390
rect 263344 1538 263504 178390
rect 271024 1538 271184 178390
rect 278704 1538 278864 178390
<< obsm4 >>
rect 5894 178420 268842 179695
rect 5894 1508 9874 178420
rect 10094 1508 17554 178420
rect 17774 1508 25234 178420
rect 25454 1508 32914 178420
rect 33134 1508 40594 178420
rect 40814 1508 48274 178420
rect 48494 1508 55954 178420
rect 56174 1508 63634 178420
rect 63854 1508 71314 178420
rect 71534 1508 78994 178420
rect 79214 1508 86674 178420
rect 86894 1508 94354 178420
rect 94574 1508 102034 178420
rect 102254 1508 109714 178420
rect 109934 1508 117394 178420
rect 117614 1508 125074 178420
rect 125294 1508 132754 178420
rect 132974 1508 140434 178420
rect 140654 1508 148114 178420
rect 148334 1508 155794 178420
rect 156014 1508 163474 178420
rect 163694 1508 171154 178420
rect 171374 1508 178834 178420
rect 179054 1508 186514 178420
rect 186734 1508 194194 178420
rect 194414 1508 201874 178420
rect 202094 1508 209554 178420
rect 209774 1508 217234 178420
rect 217454 1508 224914 178420
rect 225134 1508 232594 178420
rect 232814 1508 240274 178420
rect 240494 1508 247954 178420
rect 248174 1508 255634 178420
rect 255854 1508 263314 178420
rect 263534 1508 268842 178420
rect 5894 289 268842 1508
<< labels >>
rlabel metal2 s 174720 179600 174776 179900 6 rambus_wb_ack_o
port 1 nsew signal output
rlabel metal2 s 8400 179600 8456 179900 6 rambus_wb_addr_i[0]
port 2 nsew signal input
rlabel metal3 s 279600 107856 279900 107912 6 rambus_wb_addr_i[1]
port 3 nsew signal input
rlabel metal2 s 97104 179600 97160 179900 6 rambus_wb_addr_i[2]
port 4 nsew signal input
rlabel metal2 s 22176 100 22232 400 6 rambus_wb_addr_i[3]
port 5 nsew signal input
rlabel metal3 s 100 177408 400 177464 6 rambus_wb_addr_i[4]
port 6 nsew signal input
rlabel metal3 s 279600 41328 279900 41384 6 rambus_wb_addr_i[5]
port 7 nsew signal input
rlabel metal2 s 199584 100 199640 400 6 rambus_wb_addr_i[6]
port 8 nsew signal input
rlabel metal3 s 100 11088 400 11144 6 rambus_wb_addr_i[7]
port 9 nsew signal input
rlabel metal2 s 188496 100 188552 400 6 rambus_wb_addr_i[8]
port 10 nsew signal input
rlabel metal3 s 100 33264 400 33320 6 rambus_wb_clk_i
port 11 nsew signal input
rlabel metal3 s 100 144144 400 144200 6 rambus_wb_cyc_i
port 12 nsew signal input
rlabel metal3 s 100 55440 400 55496 6 rambus_wb_dat_i[0]
port 13 nsew signal input
rlabel metal3 s 100 133056 400 133112 6 rambus_wb_dat_i[10]
port 14 nsew signal input
rlabel metal2 s 232848 100 232904 400 6 rambus_wb_dat_i[11]
port 15 nsew signal input
rlabel metal2 s 274512 179600 274568 179900 6 rambus_wb_dat_i[12]
port 16 nsew signal input
rlabel metal2 s 41664 179600 41720 179900 6 rambus_wb_dat_i[13]
port 17 nsew signal input
rlabel metal2 s 219072 179600 219128 179900 6 rambus_wb_dat_i[14]
port 18 nsew signal input
rlabel metal2 s 266112 100 266168 400 6 rambus_wb_dat_i[15]
port 19 nsew signal input
rlabel metal2 s 163632 179600 163688 179900 6 rambus_wb_dat_i[16]
port 20 nsew signal input
rlabel metal3 s 279600 85680 279900 85736 6 rambus_wb_dat_i[17]
port 21 nsew signal input
rlabel metal3 s 279600 30240 279900 30296 6 rambus_wb_dat_i[18]
port 22 nsew signal input
rlabel metal3 s 279600 118944 279900 119000 6 rambus_wb_dat_i[19]
port 23 nsew signal input
rlabel metal2 s 30576 179600 30632 179900 6 rambus_wb_dat_i[1]
port 24 nsew signal input
rlabel metal3 s 279600 152208 279900 152264 6 rambus_wb_dat_i[20]
port 25 nsew signal input
rlabel metal2 s 119280 179600 119336 179900 6 rambus_wb_dat_i[21]
port 26 nsew signal input
rlabel metal3 s 279600 96768 279900 96824 6 rambus_wb_dat_i[22]
port 27 nsew signal input
rlabel metal3 s 279600 19152 279900 19208 6 rambus_wb_dat_i[23]
port 28 nsew signal input
rlabel metal3 s 100 44352 400 44408 6 rambus_wb_dat_i[24]
port 29 nsew signal input
rlabel metal3 s 279600 141120 279900 141176 6 rambus_wb_dat_i[25]
port 30 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 rambus_wb_dat_i[26]
port 31 nsew signal input
rlabel metal2 s 210672 100 210728 400 6 rambus_wb_dat_i[27]
port 32 nsew signal input
rlabel metal2 s 207984 179600 208040 179900 6 rambus_wb_dat_i[28]
port 33 nsew signal input
rlabel metal2 s 63840 179600 63896 179900 6 rambus_wb_dat_i[29]
port 34 nsew signal input
rlabel metal2 s 185808 179600 185864 179900 6 rambus_wb_dat_i[2]
port 35 nsew signal input
rlabel metal2 s 88704 100 88760 400 6 rambus_wb_dat_i[30]
port 36 nsew signal input
rlabel metal2 s 252336 179600 252392 179900 6 rambus_wb_dat_i[31]
port 37 nsew signal input
rlabel metal3 s 279600 130032 279900 130088 6 rambus_wb_dat_i[3]
port 38 nsew signal input
rlabel metal3 s 100 121968 400 122024 6 rambus_wb_dat_i[4]
port 39 nsew signal input
rlabel metal3 s 100 88704 400 88760 6 rambus_wb_dat_i[5]
port 40 nsew signal input
rlabel metal2 s 55440 100 55496 400 6 rambus_wb_dat_i[6]
port 41 nsew signal input
rlabel metal2 s 177408 100 177464 400 6 rambus_wb_dat_i[7]
port 42 nsew signal input
rlabel metal3 s 279600 8064 279900 8120 6 rambus_wb_dat_i[8]
port 43 nsew signal input
rlabel metal2 s 255024 100 255080 400 6 rambus_wb_dat_i[9]
port 44 nsew signal input
rlabel metal2 s 144144 100 144200 400 6 rambus_wb_dat_o[0]
port 45 nsew signal output
rlabel metal2 s 52752 179600 52808 179900 6 rambus_wb_dat_o[10]
port 46 nsew signal output
rlabel metal2 s 221760 100 221816 400 6 rambus_wb_dat_o[11]
port 47 nsew signal output
rlabel metal2 s 130368 179600 130424 179900 6 rambus_wb_dat_o[12]
port 48 nsew signal output
rlabel metal2 s 277200 100 277256 400 6 rambus_wb_dat_o[13]
port 49 nsew signal output
rlabel metal3 s 279600 52416 279900 52472 6 rambus_wb_dat_o[14]
port 50 nsew signal output
rlabel metal2 s 166320 100 166376 400 6 rambus_wb_dat_o[15]
port 51 nsew signal output
rlabel metal3 s 100 155232 400 155288 6 rambus_wb_dat_o[16]
port 52 nsew signal output
rlabel metal3 s 100 22176 400 22232 6 rambus_wb_dat_o[17]
port 53 nsew signal output
rlabel metal2 s 152544 179600 152600 179900 6 rambus_wb_dat_o[18]
port 54 nsew signal output
rlabel metal2 s 110880 100 110936 400 6 rambus_wb_dat_o[19]
port 55 nsew signal output
rlabel metal2 s 0 100 56 400 6 rambus_wb_dat_o[1]
port 56 nsew signal output
rlabel metal2 s 133056 100 133112 400 6 rambus_wb_dat_o[20]
port 57 nsew signal output
rlabel metal2 s 141456 179600 141512 179900 6 rambus_wb_dat_o[21]
port 58 nsew signal output
rlabel metal2 s 196896 179600 196952 179900 6 rambus_wb_dat_o[22]
port 59 nsew signal output
rlabel metal2 s 263424 179600 263480 179900 6 rambus_wb_dat_o[23]
port 60 nsew signal output
rlabel metal3 s 100 166320 400 166376 6 rambus_wb_dat_o[24]
port 61 nsew signal output
rlabel metal2 s 33264 100 33320 400 6 rambus_wb_dat_o[25]
port 62 nsew signal output
rlabel metal2 s 11088 100 11144 400 6 rambus_wb_dat_o[26]
port 63 nsew signal output
rlabel metal3 s 279600 174384 279900 174440 6 rambus_wb_dat_o[27]
port 64 nsew signal output
rlabel metal3 s 100 77616 400 77672 6 rambus_wb_dat_o[28]
port 65 nsew signal output
rlabel metal2 s 99792 100 99848 400 6 rambus_wb_dat_o[29]
port 66 nsew signal output
rlabel metal3 s 279600 163296 279900 163352 6 rambus_wb_dat_o[2]
port 67 nsew signal output
rlabel metal2 s 243936 100 243992 400 6 rambus_wb_dat_o[30]
port 68 nsew signal output
rlabel metal2 s 86016 179600 86072 179900 6 rambus_wb_dat_o[31]
port 69 nsew signal output
rlabel metal3 s 100 110880 400 110936 6 rambus_wb_dat_o[3]
port 70 nsew signal output
rlabel metal2 s 44352 100 44408 400 6 rambus_wb_dat_o[4]
port 71 nsew signal output
rlabel metal2 s 77616 100 77672 400 6 rambus_wb_dat_o[5]
port 72 nsew signal output
rlabel metal3 s 100 99792 400 99848 6 rambus_wb_dat_o[6]
port 73 nsew signal output
rlabel metal3 s 279600 74592 279900 74648 6 rambus_wb_dat_o[7]
port 74 nsew signal output
rlabel metal2 s 121968 100 122024 400 6 rambus_wb_dat_o[8]
port 75 nsew signal output
rlabel metal2 s 241248 179600 241304 179900 6 rambus_wb_dat_o[9]
port 76 nsew signal output
rlabel metal2 s 230160 179600 230216 179900 6 rambus_wb_rst_i
port 77 nsew signal input
rlabel metal2 s 74928 179600 74984 179900 6 rambus_wb_sel_i[0]
port 78 nsew signal input
rlabel metal2 s 108192 179600 108248 179900 6 rambus_wb_sel_i[1]
port 79 nsew signal input
rlabel metal2 s 155232 100 155288 400 6 rambus_wb_sel_i[2]
port 80 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 rambus_wb_sel_i[3]
port 81 nsew signal input
rlabel metal2 s 19488 179600 19544 179900 6 rambus_wb_stb_i
port 82 nsew signal input
rlabel metal3 s 279600 63504 279900 63560 6 rambus_wb_we_i
port 83 nsew signal input
rlabel metal4 s 2224 1538 2384 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 178390 6 vdd
port 84 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 178390 6 vss
port 85 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 178390 6 vss
port 85 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 280000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 71290680
string GDS_FILE /home/uri/p/gf180_spell/openlane/rambus/runs/22_12_05_12_50/results/signoff/rambus.magic.gds
string GDS_START 356614
<< end >>

