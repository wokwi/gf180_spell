VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spell
  CLASS BLOCK ;
  FOREIGN spell ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 896.000 27.440 899.000 ;
    END
  END clock
  PIN i_la_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1.000 803.600 4.000 ;
    END
  END i_la_addr[0]
  PIN i_la_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 661.920 4.000 662.480 ;
    END
  END i_la_addr[1]
  PIN i_la_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END i_la_addr[2]
  PIN i_la_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END i_la_addr[3]
  PIN i_la_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1.000 205.520 4.000 ;
    END
  END i_la_addr[4]
  PIN i_la_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 456.960 899.000 457.520 ;
    END
  END i_la_addr[5]
  PIN i_la_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 896.000 400.400 899.000 ;
    END
  END i_la_addr[6]
  PIN i_la_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 359.520 4.000 360.080 ;
    END
  END i_la_data[0]
  PIN i_la_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 235.200 899.000 235.760 ;
    END
  END i_la_data[1]
  PIN i_la_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END i_la_data[2]
  PIN i_la_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 719.040 4.000 719.600 ;
    END
  END i_la_data[3]
  PIN i_la_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 896.000 67.760 899.000 ;
    END
  END i_la_data[4]
  PIN i_la_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 896.000 249.200 899.000 ;
    END
  END i_la_data[5]
  PIN i_la_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 621.600 899.000 622.160 ;
    END
  END i_la_data[6]
  PIN i_la_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 896.000 649.040 899.000 ;
    END
  END i_la_data[7]
  PIN i_la_wb_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 510.720 899.000 511.280 ;
    END
  END i_la_wb_disable
  PIN i_la_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 470.400 899.000 470.960 ;
    END
  END i_la_write
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 40.320 899.000 40.880 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 1.000 218.960 4.000 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 896.000 635.600 899.000 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.320 4.000 124.880 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 896.000 622.160 899.000 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1.000 622.160 4.000 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 386.400 899.000 386.960 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.640 4.000 81.200 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 896.000 262.640 899.000 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 1.000 360.080 4.000 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 896.000 817.040 899.000 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 816.480 899.000 817.040 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.280 4.000 329.840 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.400 4.000 218.960 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 896.000 218.960 899.000 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 870.240 4.000 870.800 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 1.000 440.720 4.000 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 537.600 899.000 538.160 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1.000 733.040 4.000 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 896.000 165.200 899.000 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.640 4.000 165.200 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 1.000 40.880 4.000 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1.000 551.600 4.000 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.760 4.000 138.320 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 456.960 4.000 457.520 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 1.000 346.640 4.000 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 896.000 440.720 899.000 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 581.280 4.000 581.840 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 13.440 899.000 14.000 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 896.000 706.160 899.000 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 1.000 773.360 4.000 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 896.000 289.520 899.000 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 896.000 94.640 899.000 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1.000 497.840 4.000 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 896.000 386.960 899.000 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 896.000 0.560 899.000 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 896.000 719.600 899.000 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 678.720 899.000 679.280 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 759.360 4.000 759.920 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 359.520 899.000 360.080 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 896.000 302.960 899.000 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 896.000 870.800 899.000 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 896.000 124.880 899.000 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 483.840 899.000 484.400 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 896.000 373.520 899.000 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 164.640 899.000 165.200 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 732.480 4.000 733.040 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 275.520 899.000 276.080 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 67.200 4.000 67.760 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 0.000 899.000 0.560 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1.000 759.920 4.000 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 151.200 899.000 151.760 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 803.040 4.000 803.600 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 413.280 899.000 413.840 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.840 4.000 484.400 ;
    END
  END i_wb_data[9]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 124.320 899.000 124.880 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 719.040 899.000 719.600 ;
    END
  END i_wb_we
  PIN interrupt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 896.000 773.360 899.000 ;
    END
  END interrupt
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 843.360 4.000 843.920 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 567.840 899.000 568.400 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 1.000 817.040 4.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 896.000 470.960 899.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1.000 830.480 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 896.000 692.720 899.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 705.600 899.000 706.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 896.000 484.400 899.000 ;
    END
  END io_in[7]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 896.000 205.520 899.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 896.000 346.640 899.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 1.000 595.280 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 896.000 568.400 899.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 262.080 899.000 262.640 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 594.720 899.000 595.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END io_oeb[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 829.920 4.000 830.480 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 843.360 899.000 843.920 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.440 4.000 14.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1.000 94.640 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.600 4.000 538.160 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 896.000 497.840 899.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 896.000 413.840 899.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 896.000 40.880 899.000 ;
    END
  END io_out[7]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.320 4.000 40.880 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 896.000 897.680 899.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 896.000 759.920 899.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 896.000 524.720 899.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 635.040 4.000 635.600 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 94.080 4.000 94.640 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 896.000 457.520 899.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 1.000 706.160 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 789.600 4.000 790.160 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.280 4.000 497.840 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 772.800 4.000 773.360 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1.000 276.080 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 497.280 899.000 497.840 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 896.000 884.240 899.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 896.000 54.320 899.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1.000 484.400 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.520 4.000 276.080 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 567.840 4.000 568.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 896.000 733.040 899.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 870.240 899.000 870.800 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 896.000 360.080 899.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 107.520 899.000 108.080 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1.000 511.280 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 524.160 899.000 524.720 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 1.000 746.480 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 745.920 899.000 746.480 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1.000 635.600 4.000 ;
    END
  END la_data_out[9]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 896.000 81.200 899.000 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 896.000 276.080 899.000 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 137.760 899.000 138.320 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 248.640 899.000 249.200 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 1.000 662.480 4.000 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 470.400 4.000 470.960 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 896.000 235.760 899.000 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 346.080 899.000 346.640 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 440.160 4.000 440.720 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 896.000 803.600 899.000 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 1.000 843.920 4.000 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 67.200 899.000 67.760 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 789.600 899.000 790.160 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 896.000 857.360 899.000 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 896.000 551.600 899.000 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 524.160 4.000 524.720 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 372.960 899.000 373.520 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 329.280 899.000 329.840 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 288.960 899.000 289.520 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 80.640 899.000 81.200 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 1.000 719.600 4.000 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 856.800 899.000 857.360 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 648.480 899.000 649.040 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1.000 427.280 4.000 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 896.000 178.640 899.000 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 26.880 899.000 27.440 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 896.000 511.280 899.000 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 594.720 4.000 595.280 ;
    END
  END o_wb_data[9]
  PIN rambus_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 1.000 81.200 4.000 ;
    END
  END rambus_wb_ack_i
  PIN rambus_wb_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 896.000 662.480 899.000 ;
    END
  END rambus_wb_addr_o[0]
  PIN rambus_wb_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 346.080 4.000 346.640 ;
    END
  END rambus_wb_addr_o[1]
  PIN rambus_wb_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 608.160 899.000 608.720 ;
    END
  END rambus_wb_addr_o[2]
  PIN rambus_wb_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END rambus_wb_addr_o[3]
  PIN rambus_wb_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 803.040 899.000 803.600 ;
    END
  END rambus_wb_addr_o[4]
  PIN rambus_wb_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 204.960 899.000 205.520 ;
    END
  END rambus_wb_addr_o[5]
  PIN rambus_wb_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1.000 608.720 4.000 ;
    END
  END rambus_wb_addr_o[6]
  PIN rambus_wb_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 829.920 899.000 830.480 ;
    END
  END rambus_wb_addr_o[7]
  PIN rambus_wb_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END rambus_wb_addr_o[8]
  PIN rambus_wb_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END rambus_wb_addr_o[9]
  PIN rambus_wb_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 896.000 14.000 899.000 ;
    END
  END rambus_wb_clk_o
  PIN rambus_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1.000 790.160 4.000 ;
    END
  END rambus_wb_cyc_o
  PIN rambus_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 94.080 899.000 94.640 ;
    END
  END rambus_wb_dat_i[0]
  PIN rambus_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 896.000 581.840 899.000 ;
    END
  END rambus_wb_dat_i[10]
  PIN rambus_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 581.280 899.000 581.840 ;
    END
  END rambus_wb_dat_i[11]
  PIN rambus_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 896.000 138.320 899.000 ;
    END
  END rambus_wb_dat_i[12]
  PIN rambus_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 896.000 192.080 899.000 ;
    END
  END rambus_wb_dat_i[13]
  PIN rambus_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 896.000 151.760 899.000 ;
    END
  END rambus_wb_dat_i[14]
  PIN rambus_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END rambus_wb_dat_i[15]
  PIN rambus_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 1.000 165.200 4.000 ;
    END
  END rambus_wb_dat_i[16]
  PIN rambus_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 315.840 899.000 316.400 ;
    END
  END rambus_wb_dat_i[17]
  PIN rambus_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1.000 457.520 4.000 ;
    END
  END rambus_wb_dat_i[18]
  PIN rambus_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 896.000 830.480 899.000 ;
    END
  END rambus_wb_dat_i[19]
  PIN rambus_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 772.800 899.000 773.360 ;
    END
  END rambus_wb_dat_i[1]
  PIN rambus_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 896.000 316.400 899.000 ;
    END
  END rambus_wb_dat_i[20]
  PIN rambus_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END rambus_wb_dat_i[21]
  PIN rambus_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 399.840 899.000 400.400 ;
    END
  END rambus_wb_dat_i[22]
  PIN rambus_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 759.360 899.000 759.920 ;
    END
  END rambus_wb_dat_i[23]
  PIN rambus_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 816.480 4.000 817.040 ;
    END
  END rambus_wb_dat_i[24]
  PIN rambus_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 551.040 899.000 551.600 ;
    END
  END rambus_wb_dat_i[25]
  PIN rambus_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 191.520 899.000 192.080 ;
    END
  END rambus_wb_dat_i[26]
  PIN rambus_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 1.000 568.400 4.000 ;
    END
  END rambus_wb_dat_i[27]
  PIN rambus_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 883.680 899.000 884.240 ;
    END
  END rambus_wb_dat_i[28]
  PIN rambus_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 896.000 427.280 899.000 ;
    END
  END rambus_wb_dat_i[29]
  PIN rambus_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END rambus_wb_dat_i[2]
  PIN rambus_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 510.720 4.000 511.280 ;
    END
  END rambus_wb_dat_i[30]
  PIN rambus_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 372.960 4.000 373.520 ;
    END
  END rambus_wb_dat_i[31]
  PIN rambus_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 178.080 899.000 178.640 ;
    END
  END rambus_wb_dat_i[3]
  PIN rambus_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 705.600 4.000 706.160 ;
    END
  END rambus_wb_dat_i[4]
  PIN rambus_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 1.000 870.800 4.000 ;
    END
  END rambus_wb_dat_i[5]
  PIN rambus_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 1.000 138.320 4.000 ;
    END
  END rambus_wb_dat_i[6]
  PIN rambus_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END rambus_wb_dat_i[7]
  PIN rambus_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 302.400 899.000 302.960 ;
    END
  END rambus_wb_dat_i[8]
  PIN rambus_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 896.000 843.920 899.000 ;
    END
  END rambus_wb_dat_i[9]
  PIN rambus_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 692.160 899.000 692.720 ;
    END
  END rambus_wb_dat_o[0]
  PIN rambus_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 1.000 884.240 4.000 ;
    END
  END rambus_wb_dat_o[10]
  PIN rambus_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 1.000 67.760 4.000 ;
    END
  END rambus_wb_dat_o[11]
  PIN rambus_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 426.720 899.000 427.280 ;
    END
  END rambus_wb_dat_o[12]
  PIN rambus_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1.000 14.000 4.000 ;
    END
  END rambus_wb_dat_o[13]
  PIN rambus_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 732.480 899.000 733.040 ;
    END
  END rambus_wb_dat_o[14]
  PIN rambus_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 896.000 790.160 899.000 ;
    END
  END rambus_wb_dat_o[15]
  PIN rambus_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 53.760 899.000 54.320 ;
    END
  END rambus_wb_dat_o[16]
  PIN rambus_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 896.000 746.480 899.000 ;
    END
  END rambus_wb_dat_o[17]
  PIN rambus_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END rambus_wb_dat_o[18]
  PIN rambus_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.720 4.000 427.280 ;
    END
  END rambus_wb_dat_o[19]
  PIN rambus_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 1.000 581.840 4.000 ;
    END
  END rambus_wb_dat_o[1]
  PIN rambus_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END rambus_wb_dat_o[20]
  PIN rambus_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END rambus_wb_dat_o[21]
  PIN rambus_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 551.040 4.000 551.600 ;
    END
  END rambus_wb_dat_o[22]
  PIN rambus_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 883.680 4.000 884.240 ;
    END
  END rambus_wb_dat_o[23]
  PIN rambus_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END rambus_wb_dat_o[24]
  PIN rambus_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END rambus_wb_dat_o[25]
  PIN rambus_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END rambus_wb_dat_o[26]
  PIN rambus_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END rambus_wb_dat_o[27]
  PIN rambus_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 896.000 538.160 899.000 ;
    END
  END rambus_wb_dat_o[28]
  PIN rambus_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 896.000 329.840 899.000 ;
    END
  END rambus_wb_dat_o[29]
  PIN rambus_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 1.000 470.960 4.000 ;
    END
  END rambus_wb_dat_o[2]
  PIN rambus_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 896.000 679.280 899.000 ;
    END
  END rambus_wb_dat_o[30]
  PIN rambus_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 218.400 899.000 218.960 ;
    END
  END rambus_wb_dat_o[31]
  PIN rambus_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 648.480 4.000 649.040 ;
    END
  END rambus_wb_dat_o[3]
  PIN rambus_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 661.920 899.000 662.480 ;
    END
  END rambus_wb_dat_o[4]
  PIN rambus_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END rambus_wb_dat_o[5]
  PIN rambus_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1.000 329.840 4.000 ;
    END
  END rambus_wb_dat_o[6]
  PIN rambus_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 1.000 524.720 4.000 ;
    END
  END rambus_wb_dat_o[7]
  PIN rambus_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 635.040 899.000 635.600 ;
    END
  END rambus_wb_dat_o[8]
  PIN rambus_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1.000 538.160 4.000 ;
    END
  END rambus_wb_dat_o[9]
  PIN rambus_wb_rst_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 896.000 608.720 899.000 ;
    END
  END rambus_wb_rst_o
  PIN rambus_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 896.000 595.280 899.000 ;
    END
  END rambus_wb_sel_o[0]
  PIN rambus_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END rambus_wb_sel_o[1]
  PIN rambus_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 896.000 108.080 899.000 ;
    END
  END rambus_wb_sel_o[2]
  PIN rambus_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 1.000 649.040 4.000 ;
    END
  END rambus_wb_sel_o[3]
  PIN rambus_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.960 4.000 205.520 ;
    END
  END rambus_wb_stb_o
  PIN rambus_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 745.920 4.000 746.480 ;
    END
  END rambus_wb_we_o
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 896.000 440.160 899.000 440.720 ;
    END
  END reset
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 882.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 882.300 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 893.200 882.300 ;
      LAYER Metal2 ;
        RECT 0.860 895.700 13.140 896.000 ;
        RECT 14.300 895.700 26.580 896.000 ;
        RECT 27.740 895.700 40.020 896.000 ;
        RECT 41.180 895.700 53.460 896.000 ;
        RECT 54.620 895.700 66.900 896.000 ;
        RECT 68.060 895.700 80.340 896.000 ;
        RECT 81.500 895.700 93.780 896.000 ;
        RECT 94.940 895.700 107.220 896.000 ;
        RECT 108.380 895.700 124.020 896.000 ;
        RECT 125.180 895.700 137.460 896.000 ;
        RECT 138.620 895.700 150.900 896.000 ;
        RECT 152.060 895.700 164.340 896.000 ;
        RECT 165.500 895.700 177.780 896.000 ;
        RECT 178.940 895.700 191.220 896.000 ;
        RECT 192.380 895.700 204.660 896.000 ;
        RECT 205.820 895.700 218.100 896.000 ;
        RECT 219.260 895.700 234.900 896.000 ;
        RECT 236.060 895.700 248.340 896.000 ;
        RECT 249.500 895.700 261.780 896.000 ;
        RECT 262.940 895.700 275.220 896.000 ;
        RECT 276.380 895.700 288.660 896.000 ;
        RECT 289.820 895.700 302.100 896.000 ;
        RECT 303.260 895.700 315.540 896.000 ;
        RECT 316.700 895.700 328.980 896.000 ;
        RECT 330.140 895.700 345.780 896.000 ;
        RECT 346.940 895.700 359.220 896.000 ;
        RECT 360.380 895.700 372.660 896.000 ;
        RECT 373.820 895.700 386.100 896.000 ;
        RECT 387.260 895.700 399.540 896.000 ;
        RECT 400.700 895.700 412.980 896.000 ;
        RECT 414.140 895.700 426.420 896.000 ;
        RECT 427.580 895.700 439.860 896.000 ;
        RECT 441.020 895.700 456.660 896.000 ;
        RECT 457.820 895.700 470.100 896.000 ;
        RECT 471.260 895.700 483.540 896.000 ;
        RECT 484.700 895.700 496.980 896.000 ;
        RECT 498.140 895.700 510.420 896.000 ;
        RECT 511.580 895.700 523.860 896.000 ;
        RECT 525.020 895.700 537.300 896.000 ;
        RECT 538.460 895.700 550.740 896.000 ;
        RECT 551.900 895.700 567.540 896.000 ;
        RECT 568.700 895.700 580.980 896.000 ;
        RECT 582.140 895.700 594.420 896.000 ;
        RECT 595.580 895.700 607.860 896.000 ;
        RECT 609.020 895.700 621.300 896.000 ;
        RECT 622.460 895.700 634.740 896.000 ;
        RECT 635.900 895.700 648.180 896.000 ;
        RECT 649.340 895.700 661.620 896.000 ;
        RECT 662.780 895.700 678.420 896.000 ;
        RECT 679.580 895.700 691.860 896.000 ;
        RECT 693.020 895.700 705.300 896.000 ;
        RECT 706.460 895.700 718.740 896.000 ;
        RECT 719.900 895.700 732.180 896.000 ;
        RECT 733.340 895.700 745.620 896.000 ;
        RECT 746.780 895.700 759.060 896.000 ;
        RECT 760.220 895.700 772.500 896.000 ;
        RECT 773.660 895.700 789.300 896.000 ;
        RECT 790.460 895.700 802.740 896.000 ;
        RECT 803.900 895.700 816.180 896.000 ;
        RECT 817.340 895.700 829.620 896.000 ;
        RECT 830.780 895.700 843.060 896.000 ;
        RECT 844.220 895.700 856.500 896.000 ;
        RECT 857.660 895.700 869.940 896.000 ;
        RECT 871.100 895.700 883.380 896.000 ;
        RECT 884.540 895.700 896.820 896.000 ;
        RECT 0.140 4.300 897.540 895.700 ;
        RECT 0.860 0.700 13.140 4.300 ;
        RECT 14.300 0.700 26.580 4.300 ;
        RECT 27.740 0.700 40.020 4.300 ;
        RECT 41.180 0.700 53.460 4.300 ;
        RECT 54.620 0.700 66.900 4.300 ;
        RECT 68.060 0.700 80.340 4.300 ;
        RECT 81.500 0.700 93.780 4.300 ;
        RECT 94.940 0.700 107.220 4.300 ;
        RECT 108.380 0.700 124.020 4.300 ;
        RECT 125.180 0.700 137.460 4.300 ;
        RECT 138.620 0.700 150.900 4.300 ;
        RECT 152.060 0.700 164.340 4.300 ;
        RECT 165.500 0.700 177.780 4.300 ;
        RECT 178.940 0.700 191.220 4.300 ;
        RECT 192.380 0.700 204.660 4.300 ;
        RECT 205.820 0.700 218.100 4.300 ;
        RECT 219.260 0.700 234.900 4.300 ;
        RECT 236.060 0.700 248.340 4.300 ;
        RECT 249.500 0.700 261.780 4.300 ;
        RECT 262.940 0.700 275.220 4.300 ;
        RECT 276.380 0.700 288.660 4.300 ;
        RECT 289.820 0.700 302.100 4.300 ;
        RECT 303.260 0.700 315.540 4.300 ;
        RECT 316.700 0.700 328.980 4.300 ;
        RECT 330.140 0.700 345.780 4.300 ;
        RECT 346.940 0.700 359.220 4.300 ;
        RECT 360.380 0.700 372.660 4.300 ;
        RECT 373.820 0.700 386.100 4.300 ;
        RECT 387.260 0.700 399.540 4.300 ;
        RECT 400.700 0.700 412.980 4.300 ;
        RECT 414.140 0.700 426.420 4.300 ;
        RECT 427.580 0.700 439.860 4.300 ;
        RECT 441.020 0.700 456.660 4.300 ;
        RECT 457.820 0.700 470.100 4.300 ;
        RECT 471.260 0.700 483.540 4.300 ;
        RECT 484.700 0.700 496.980 4.300 ;
        RECT 498.140 0.700 510.420 4.300 ;
        RECT 511.580 0.700 523.860 4.300 ;
        RECT 525.020 0.700 537.300 4.300 ;
        RECT 538.460 0.700 550.740 4.300 ;
        RECT 551.900 0.700 567.540 4.300 ;
        RECT 568.700 0.700 580.980 4.300 ;
        RECT 582.140 0.700 594.420 4.300 ;
        RECT 595.580 0.700 607.860 4.300 ;
        RECT 609.020 0.700 621.300 4.300 ;
        RECT 622.460 0.700 634.740 4.300 ;
        RECT 635.900 0.700 648.180 4.300 ;
        RECT 649.340 0.700 661.620 4.300 ;
        RECT 662.780 0.700 678.420 4.300 ;
        RECT 679.580 0.700 691.860 4.300 ;
        RECT 693.020 0.700 705.300 4.300 ;
        RECT 706.460 0.700 718.740 4.300 ;
        RECT 719.900 0.700 732.180 4.300 ;
        RECT 733.340 0.700 745.620 4.300 ;
        RECT 746.780 0.700 759.060 4.300 ;
        RECT 760.220 0.700 772.500 4.300 ;
        RECT 773.660 0.700 789.300 4.300 ;
        RECT 790.460 0.700 802.740 4.300 ;
        RECT 803.900 0.700 816.180 4.300 ;
        RECT 817.340 0.700 829.620 4.300 ;
        RECT 830.780 0.700 843.060 4.300 ;
        RECT 844.220 0.700 856.500 4.300 ;
        RECT 857.660 0.700 869.940 4.300 ;
        RECT 871.100 0.700 883.380 4.300 ;
        RECT 884.540 0.700 897.540 4.300 ;
        RECT 0.140 0.090 897.540 0.700 ;
      LAYER Metal3 ;
        RECT 0.090 884.540 897.590 890.820 ;
        RECT 0.090 883.380 0.700 884.540 ;
        RECT 4.300 883.380 895.700 884.540 ;
        RECT 0.090 871.100 897.590 883.380 ;
        RECT 0.090 869.940 0.700 871.100 ;
        RECT 4.300 869.940 895.700 871.100 ;
        RECT 0.090 857.660 897.590 869.940 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 895.700 857.660 ;
        RECT 0.090 844.220 897.590 856.500 ;
        RECT 0.090 843.060 0.700 844.220 ;
        RECT 4.300 843.060 895.700 844.220 ;
        RECT 0.090 830.780 897.590 843.060 ;
        RECT 0.090 829.620 0.700 830.780 ;
        RECT 4.300 829.620 895.700 830.780 ;
        RECT 0.090 817.340 897.590 829.620 ;
        RECT 0.090 816.180 0.700 817.340 ;
        RECT 4.300 816.180 895.700 817.340 ;
        RECT 0.090 803.900 897.590 816.180 ;
        RECT 0.090 802.740 0.700 803.900 ;
        RECT 4.300 802.740 895.700 803.900 ;
        RECT 0.090 790.460 897.590 802.740 ;
        RECT 0.090 789.300 0.700 790.460 ;
        RECT 4.300 789.300 895.700 790.460 ;
        RECT 0.090 773.660 897.590 789.300 ;
        RECT 0.090 772.500 0.700 773.660 ;
        RECT 4.300 772.500 895.700 773.660 ;
        RECT 0.090 760.220 897.590 772.500 ;
        RECT 0.090 759.060 0.700 760.220 ;
        RECT 4.300 759.060 895.700 760.220 ;
        RECT 0.090 746.780 897.590 759.060 ;
        RECT 0.090 745.620 0.700 746.780 ;
        RECT 4.300 745.620 895.700 746.780 ;
        RECT 0.090 733.340 897.590 745.620 ;
        RECT 0.090 732.180 0.700 733.340 ;
        RECT 4.300 732.180 895.700 733.340 ;
        RECT 0.090 719.900 897.590 732.180 ;
        RECT 0.090 718.740 0.700 719.900 ;
        RECT 4.300 718.740 895.700 719.900 ;
        RECT 0.090 706.460 897.590 718.740 ;
        RECT 0.090 705.300 0.700 706.460 ;
        RECT 4.300 705.300 895.700 706.460 ;
        RECT 0.090 693.020 897.590 705.300 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 895.700 693.020 ;
        RECT 0.090 679.580 897.590 691.860 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 895.700 679.580 ;
        RECT 0.090 662.780 897.590 678.420 ;
        RECT 0.090 661.620 0.700 662.780 ;
        RECT 4.300 661.620 895.700 662.780 ;
        RECT 0.090 649.340 897.590 661.620 ;
        RECT 0.090 648.180 0.700 649.340 ;
        RECT 4.300 648.180 895.700 649.340 ;
        RECT 0.090 635.900 897.590 648.180 ;
        RECT 0.090 634.740 0.700 635.900 ;
        RECT 4.300 634.740 895.700 635.900 ;
        RECT 0.090 622.460 897.590 634.740 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 895.700 622.460 ;
        RECT 0.090 609.020 897.590 621.300 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 895.700 609.020 ;
        RECT 0.090 595.580 897.590 607.860 ;
        RECT 0.090 594.420 0.700 595.580 ;
        RECT 4.300 594.420 895.700 595.580 ;
        RECT 0.090 582.140 897.590 594.420 ;
        RECT 0.090 580.980 0.700 582.140 ;
        RECT 4.300 580.980 895.700 582.140 ;
        RECT 0.090 568.700 897.590 580.980 ;
        RECT 0.090 567.540 0.700 568.700 ;
        RECT 4.300 567.540 895.700 568.700 ;
        RECT 0.090 551.900 897.590 567.540 ;
        RECT 0.090 550.740 0.700 551.900 ;
        RECT 4.300 550.740 895.700 551.900 ;
        RECT 0.090 538.460 897.590 550.740 ;
        RECT 0.090 537.300 0.700 538.460 ;
        RECT 4.300 537.300 895.700 538.460 ;
        RECT 0.090 525.020 897.590 537.300 ;
        RECT 0.090 523.860 0.700 525.020 ;
        RECT 4.300 523.860 895.700 525.020 ;
        RECT 0.090 511.580 897.590 523.860 ;
        RECT 0.090 510.420 0.700 511.580 ;
        RECT 4.300 510.420 895.700 511.580 ;
        RECT 0.090 498.140 897.590 510.420 ;
        RECT 0.090 496.980 0.700 498.140 ;
        RECT 4.300 496.980 895.700 498.140 ;
        RECT 0.090 484.700 897.590 496.980 ;
        RECT 0.090 483.540 0.700 484.700 ;
        RECT 4.300 483.540 895.700 484.700 ;
        RECT 0.090 471.260 897.590 483.540 ;
        RECT 0.090 470.100 0.700 471.260 ;
        RECT 4.300 470.100 895.700 471.260 ;
        RECT 0.090 457.820 897.590 470.100 ;
        RECT 0.090 456.660 0.700 457.820 ;
        RECT 4.300 456.660 895.700 457.820 ;
        RECT 0.090 441.020 897.590 456.660 ;
        RECT 0.090 439.860 0.700 441.020 ;
        RECT 4.300 439.860 895.700 441.020 ;
        RECT 0.090 427.580 897.590 439.860 ;
        RECT 0.090 426.420 0.700 427.580 ;
        RECT 4.300 426.420 895.700 427.580 ;
        RECT 0.090 414.140 897.590 426.420 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 895.700 414.140 ;
        RECT 0.090 400.700 897.590 412.980 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 895.700 400.700 ;
        RECT 0.090 387.260 897.590 399.540 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 895.700 387.260 ;
        RECT 0.090 373.820 897.590 386.100 ;
        RECT 0.090 372.660 0.700 373.820 ;
        RECT 4.300 372.660 895.700 373.820 ;
        RECT 0.090 360.380 897.590 372.660 ;
        RECT 0.090 359.220 0.700 360.380 ;
        RECT 4.300 359.220 895.700 360.380 ;
        RECT 0.090 346.940 897.590 359.220 ;
        RECT 0.090 345.780 0.700 346.940 ;
        RECT 4.300 345.780 895.700 346.940 ;
        RECT 0.090 330.140 897.590 345.780 ;
        RECT 0.090 328.980 0.700 330.140 ;
        RECT 4.300 328.980 895.700 330.140 ;
        RECT 0.090 316.700 897.590 328.980 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 895.700 316.700 ;
        RECT 0.090 303.260 897.590 315.540 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 895.700 303.260 ;
        RECT 0.090 289.820 897.590 302.100 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 895.700 289.820 ;
        RECT 0.090 276.380 897.590 288.660 ;
        RECT 0.090 275.220 0.700 276.380 ;
        RECT 4.300 275.220 895.700 276.380 ;
        RECT 0.090 262.940 897.590 275.220 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 895.700 262.940 ;
        RECT 0.090 249.500 897.590 261.780 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 895.700 249.500 ;
        RECT 0.090 236.060 897.590 248.340 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 895.700 236.060 ;
        RECT 0.090 219.260 897.590 234.900 ;
        RECT 0.090 218.100 0.700 219.260 ;
        RECT 4.300 218.100 895.700 219.260 ;
        RECT 0.090 205.820 897.590 218.100 ;
        RECT 0.090 204.660 0.700 205.820 ;
        RECT 4.300 204.660 895.700 205.820 ;
        RECT 0.090 192.380 897.590 204.660 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 895.700 192.380 ;
        RECT 0.090 178.940 897.590 191.220 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 895.700 178.940 ;
        RECT 0.090 165.500 897.590 177.780 ;
        RECT 0.090 164.340 0.700 165.500 ;
        RECT 4.300 164.340 895.700 165.500 ;
        RECT 0.090 152.060 897.590 164.340 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 895.700 152.060 ;
        RECT 0.090 138.620 897.590 150.900 ;
        RECT 0.090 137.460 0.700 138.620 ;
        RECT 4.300 137.460 895.700 138.620 ;
        RECT 0.090 125.180 897.590 137.460 ;
        RECT 0.090 124.020 0.700 125.180 ;
        RECT 4.300 124.020 895.700 125.180 ;
        RECT 0.090 108.380 897.590 124.020 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 895.700 108.380 ;
        RECT 0.090 94.940 897.590 107.220 ;
        RECT 0.090 93.780 0.700 94.940 ;
        RECT 4.300 93.780 895.700 94.940 ;
        RECT 0.090 81.500 897.590 93.780 ;
        RECT 0.090 80.340 0.700 81.500 ;
        RECT 4.300 80.340 895.700 81.500 ;
        RECT 0.090 68.060 897.590 80.340 ;
        RECT 0.090 66.900 0.700 68.060 ;
        RECT 4.300 66.900 895.700 68.060 ;
        RECT 0.090 54.620 897.590 66.900 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 895.700 54.620 ;
        RECT 0.090 41.180 897.590 53.460 ;
        RECT 0.090 40.020 0.700 41.180 ;
        RECT 4.300 40.020 895.700 41.180 ;
        RECT 0.090 27.740 897.590 40.020 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 895.700 27.740 ;
        RECT 0.090 14.300 897.590 26.580 ;
        RECT 0.090 13.140 0.700 14.300 ;
        RECT 4.300 13.140 895.700 14.300 ;
        RECT 0.090 0.860 897.590 13.140 ;
        RECT 0.090 0.140 895.700 0.860 ;
      LAYER Metal4 ;
        RECT 198.380 15.080 252.340 875.190 ;
        RECT 254.540 15.080 329.140 875.190 ;
        RECT 331.340 15.080 405.940 875.190 ;
        RECT 408.140 15.080 482.740 875.190 ;
        RECT 484.940 15.080 559.540 875.190 ;
        RECT 561.740 15.080 636.340 875.190 ;
        RECT 638.540 15.080 713.140 875.190 ;
        RECT 715.340 15.080 726.740 875.190 ;
        RECT 198.380 4.570 726.740 15.080 ;
  END
END spell
END LIBRARY

