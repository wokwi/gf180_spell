* NGSPICE file created from spell.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

.subckt spell clock i_la_addr[0] i_la_addr[1] i_la_addr[2] i_la_addr[3] i_la_addr[4]
+ i_la_addr[5] i_la_addr[6] i_la_data[0] i_la_data[1] i_la_data[2] i_la_data[3] i_la_data[4]
+ i_la_data[5] i_la_data[6] i_la_data[7] i_la_wb_disable i_la_write i_wb_addr[0] i_wb_addr[10]
+ i_wb_addr[11] i_wb_addr[12] i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16]
+ i_wb_addr[17] i_wb_addr[18] i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21]
+ i_wb_addr[22] i_wb_addr[23] i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27]
+ i_wb_addr[28] i_wb_addr[29] i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3]
+ i_wb_addr[4] i_wb_addr[5] i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc
+ i_wb_data[0] i_wb_data[10] i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14]
+ i_wb_data[15] i_wb_data[16] i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1]
+ i_wb_data[20] i_wb_data[21] i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25]
+ i_wb_data[26] i_wb_data[27] i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30]
+ i_wb_data[31] i_wb_data[3] i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8]
+ i_wb_data[9] i_wb_stb i_wb_we interrupt io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3]
+ la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ o_wb_ack o_wb_data[0] o_wb_data[10] o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14]
+ o_wb_data[15] o_wb_data[16] o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1]
+ o_wb_data[20] o_wb_data[21] o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25]
+ o_wb_data[26] o_wb_data[27] o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30]
+ o_wb_data[31] o_wb_data[3] o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8]
+ o_wb_data[9] rambus_wb_ack_i rambus_wb_addr_o[0] rambus_wb_addr_o[1] rambus_wb_addr_o[2]
+ rambus_wb_addr_o[3] rambus_wb_addr_o[4] rambus_wb_addr_o[5] rambus_wb_addr_o[6]
+ rambus_wb_addr_o[7] rambus_wb_addr_o[8] rambus_wb_addr_o[9] rambus_wb_clk_o rambus_wb_cyc_o
+ rambus_wb_dat_i[0] rambus_wb_dat_i[10] rambus_wb_dat_i[11] rambus_wb_dat_i[12] rambus_wb_dat_i[13]
+ rambus_wb_dat_i[14] rambus_wb_dat_i[15] rambus_wb_dat_i[16] rambus_wb_dat_i[17]
+ rambus_wb_dat_i[18] rambus_wb_dat_i[19] rambus_wb_dat_i[1] rambus_wb_dat_i[20] rambus_wb_dat_i[21]
+ rambus_wb_dat_i[22] rambus_wb_dat_i[23] rambus_wb_dat_i[24] rambus_wb_dat_i[25]
+ rambus_wb_dat_i[26] rambus_wb_dat_i[27] rambus_wb_dat_i[28] rambus_wb_dat_i[29]
+ rambus_wb_dat_i[2] rambus_wb_dat_i[30] rambus_wb_dat_i[31] rambus_wb_dat_i[3] rambus_wb_dat_i[4]
+ rambus_wb_dat_i[5] rambus_wb_dat_i[6] rambus_wb_dat_i[7] rambus_wb_dat_i[8] rambus_wb_dat_i[9]
+ rambus_wb_dat_o[0] rambus_wb_dat_o[10] rambus_wb_dat_o[11] rambus_wb_dat_o[12] rambus_wb_dat_o[13]
+ rambus_wb_dat_o[14] rambus_wb_dat_o[15] rambus_wb_dat_o[16] rambus_wb_dat_o[17]
+ rambus_wb_dat_o[18] rambus_wb_dat_o[19] rambus_wb_dat_o[1] rambus_wb_dat_o[20] rambus_wb_dat_o[21]
+ rambus_wb_dat_o[22] rambus_wb_dat_o[23] rambus_wb_dat_o[24] rambus_wb_dat_o[25]
+ rambus_wb_dat_o[26] rambus_wb_dat_o[27] rambus_wb_dat_o[28] rambus_wb_dat_o[29]
+ rambus_wb_dat_o[2] rambus_wb_dat_o[30] rambus_wb_dat_o[31] rambus_wb_dat_o[3] rambus_wb_dat_o[4]
+ rambus_wb_dat_o[5] rambus_wb_dat_o[6] rambus_wb_dat_o[7] rambus_wb_dat_o[8] rambus_wb_dat_o[9]
+ rambus_wb_rst_o rambus_wb_sel_o[0] rambus_wb_sel_o[1] rambus_wb_sel_o[2] rambus_wb_sel_o[3]
+ rambus_wb_stb_o rambus_wb_we_o reset vdd vss
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05903_ _01437_ _01445_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06883_ _02246_ _02335_ _02331_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09671_ _04591_ _04601_ _04628_ _04630_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07534__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05834_ _01291_ _01373_ _01377_ _01306_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08622_ _03762_ _03742_ _03763_ net148 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05832__S _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05765_ stack\[24\]\[2\] stack\[25\]\[2\] _00901_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08553_ _03703_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07504_ _02823_ _02817_ _02825_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08484_ _03217_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input108_I rambus_wb_dat_i[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05696_ _01239_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _02726_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09039__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__B2 stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07366_ _02702_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06317_ _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09105_ _03731_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07297_ _02604_ _02664_ _02660_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10417__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09036_ _04013_ _04069_ _04078_ stack\[9\]\[5\] _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input73_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06462__I _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06248_ _01211_ _01737_ _01778_ _01789_ _01719_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_164_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _01721_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06025__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06025__B2 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10567__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09938_ _04829_ _04837_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09869_ _04540_ _04785_ _04780_ net49 _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06328__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__B1 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05536__B1 stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06637__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10713_ _00305_ clknet_leaf_29_clock mem.mem_dff.data_mem\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05839__B2 _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _00236_ clknet_leaf_119_clock mem.mem_dff.code_mem\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ _00167_ clknet_leaf_89_clock mem.mem_dff.code_mem\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06264__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05311__I0 stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09202__A1 _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A2 _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07764__A1 _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11127_ _00719_ clknet_leaf_156_clock stack\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_142_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05716__I _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _00650_ clknet_leaf_22_clock delay_cycles\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09505__A2 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06319__A2 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10009_ _04881_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05550_ stack\[7\]\[6\] _01062_ _01098_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07819__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05481_ _00928_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08492__A2 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _02365_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09858__I _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07151_ _02485_ _02550_ _02546_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09441__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07378__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06102_ _01575_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07082_ _02494_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06033_ _01193_ _01234_ _01219_ _01235_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06007__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06007__B2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _01597_ _01606_ _01615_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06231__B _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05626__I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09723_ _04256_ _04659_ _04682_ _02010_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06935_ _02375_ _02364_ _02379_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07507__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _04610_ _04611_ _04564_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08937__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06866_ _02317_ _02323_ _02325_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _03747_ _03750_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05817_ stack\[18\]\[7\] stack\[19\]\[7\] _01360_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06797_ _02251_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09585_ delay_cycles\[10\] _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05748_ _01267_ _01288_ _01289_ _01291_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08536_ _03691_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05679_ _01222_ net133 net132 net131 _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_23_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08467_ _01684_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06494__A1 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05297__A2 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ mem.mem_dff.code_mem\[24\]\[0\] _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10290__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08398_ net122 _03573_ _03576_ _03079_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _02702_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09432__A1 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06246__A1 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10360_ _05156_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07994__A1 stack\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05844__I1 stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ _03827_ _03993_ _03944_ _03675_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_10291_ _03740_ _05109_ _05110_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09196__B1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09008__I _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A1 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06021__I1 stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05780__I0 stack\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08474__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10281__A2 _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10732__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _00219_ clknet_leaf_101_clock mem.mem_dff.code_mem\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09423__A1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10033__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10558_ _00150_ clknet_leaf_91_clock mem.mem_dff.code_mem\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07985__A1 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10489_ _00081_ clknet_leaf_118_clock mem.mem_dff.code_mem\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10882__CLK clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06986__B _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06720_ mem.mem_dff.code_mem\[5\]\[3\] _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08757__I _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__A1 mem.mem_dff.code_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06651_ _02138_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05602_ _01084_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ _02097_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09370_ net107 _03099_ _02618_ net102 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08321_ mem.dff_data_out\[5\] _03511_ _03483_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05533_ _01076_ _01079_ _01081_ _01040_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ mem.mem_dff.data_mem\[1\]\[3\] _03377_ _03378_ mem.mem_dff.data_mem\[3\]\[3\]
+ mem.mem_dff.data_mem\[7\]\[3\] _03379_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_178_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05464_ _01014_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10272__A2 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07203_ _02350_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03069_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08217__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09414__A1 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05395_ stack\[7\]\[3\] _00905_ _00943_ _00946_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ _02537_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06779__A2 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ _02394_ _02473_ _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05826__I1 stack\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput220 net220 rambus_wb_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07836__I mem.mem_dff.data_mem\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput231 net231 rambus_wb_stb_o vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06016_ stack\[4\]\[1\] stack\[5\]\[1\] _01472_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07728__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10262__I _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07057__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I i_wb_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07967_ _03005_ _03178_ _03181_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06951__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _04250_ _04251_ _04256_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06918_ _02365_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07898_ _03132_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08153__A1 mem.mem_dff.code_mem\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09637_ cycles_per_ms\[1\] _04596_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06849_ mem.mem_dff.code_mem\[8\]\[6\] _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__I3 stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09568_ _04513_ _04518_ _04523_ _04527_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_43_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10755__CLK clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03185_ _03676_ _03680_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _01661_ _01694_ _01257_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10263__A2 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__A1 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10412_ _00004_ clknet_leaf_169_clock stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05690__A2 _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A1 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05817__I1 stack\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _05068_ _05138_ _05145_ stack\[16\]\[6\] _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09169__B1 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06650__I _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09708__A2 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10274_ _01825_ _05090_ _05095_ stack\[30\]\[2\] _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08392__A1 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_15_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_181_clock clknet_4_4_0_clock clknet_leaf_181_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07481__I mem.mem_dff.code_mem\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A1 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10121__B _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08695__A2 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05930__S _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09644__A1 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06825__I _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08245__C _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05681__A2 _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134_clock clknet_4_6_0_clock clknet_leaf_134_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06630__A1 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06560__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__I _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _01828_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10628__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09871__I _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08383__A1 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07821_ _02030_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_149_clock clknet_4_5_0_clock clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_215_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__A1 cycles_per_ms\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07752_ _03019_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08487__I _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A1 _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06703_ _02165_ _02187_ _02195_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10778__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__S _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07683_ mem.mem_dff.code_mem\[31\]\[2\] _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09883__A1 cycles_per_ms\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08686__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__B2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__I3 stack\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09422_ _04395_ _04389_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06634_ _02132_ _02139_ _02141_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05744__I0 stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05840__S _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _04320_ _04331_ _04332_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06565_ _02072_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ _03489_ _03492_ _03493_ _03494_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10245__A2 _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05516_ stack\[14\]\[5\] _01045_ _01064_ _01065_ _00961_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06496_ _02018_ _02027_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09284_ net78 _02289_ _00760_ net94 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ _02257_ _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05447_ _00937_ _00997_ _00879_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_197_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08166_ _03351_ _03354_ _03357_ _03360_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05378_ _00925_ _00929_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07949__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07117_ _02522_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05795__B _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08097_ _02700_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08610__A2 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07566__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07048_ _02288_ _02319_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06470__I _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09781__I _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output142_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _04006_ _04048_ _04046_ stack\[25\]\[2\] _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_189_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 mem.mem_dff.data_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09323__B1 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10961_ _00553_ clknet_leaf_149_clock stack\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09874__A1 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09874__B2 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10892_ _00484_ clknet_leaf_0_clock stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05360__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06645__I _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__I _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09956__I _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_51_clock clknet_4_11_0_clock clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08860__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11083__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__A2 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06612__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__A2 _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10326_ _05133_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_clock clknet_4_11_0_clock clknet_leaf_66_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10257_ stack\[14\]\[6\] _05078_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08365__A1 mem.mem_dff.code_mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05925__S _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10188_ net173 _05035_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__A1 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10920__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05274__S1 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__I0 stack\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08668__A2 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06350_ stack\[2\]\[4\] _01830_ _01888_ _01714_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09093__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05301_ _00768_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ _01228_ _01820_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__A2 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_19_clock clknet_4_8_0_clock clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_200_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05232_ _00784_ _00785_ _00786_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08020_ _01921_ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05654__A2 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10450__CLK clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07386__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05257__I2 stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ delay_cycles\[20\] _04854_ _04859_ _04626_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _03678_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08356__A1 mem.mem_dff.code_mem\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08853_ _03942_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10163__A1 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05709__A3 _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ _03056_ _03057_ _03059_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_190_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08784_ _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05965__I0 stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08108__A1 _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05996_ _01467_ _01538_ _01539_ _01434_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07735_ mem.mem_dff.data_mem\[0\]\[5\] _03003_ _02999_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05590__A1 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__A1 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08659__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__B2 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ mem.mem_dff.code_mem\[30\]\[7\] _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09405_ _01762_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06617_ mem.mem_dff.code_mem\[2\]\[7\] _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07597_ _02897_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09336_ net90 _03042_ _03014_ net81 _04306_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05893__A2 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06465__I _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06548_ _02018_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_205_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09084__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09267_ net141 _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06479_ _02006_ _02011_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08831__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ mem.mem_dff.code_mem\[0\]\[2\] _03290_ _03401_ _03411_ _03316_ _03412_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_126_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__I _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09198_ _04131_ _04186_ _04200_ stack\[20\]\[5\] _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08149_ _02761_ _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06414__B _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ _00752_ clknet_leaf_167_clock stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10111_ _04955_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10943__CLK clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__I3 stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11091_ _00683_ clknet_leaf_14_clock net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05745__S _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04903_ _04904_ _04908_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08898__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09016__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05544__I _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09847__A1 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10944_ _00536_ clknet_leaf_142_clock stack\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _00467_ clknet_leaf_192_clock stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A2 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07086__A1 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__I _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08035__B1 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08586__A1 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09783__B1 _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10309_ stack\[27\]\[4\] _05118_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10145__A1 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08889__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05850_ _01271_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05947__I0 stack\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05781_ _01011_ _01323_ _01324_ _01286_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05572__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07520_ _02752_ _02832_ _02827_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07313__A2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11191__I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06402_ _01936_ _01938_ _01901_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10816__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07382_ _02255_ _02586_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _04145_ _04025_ _04026_ _01712_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06333_ _01866_ _01871_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08274__B1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08813__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05627__A2 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09052_ _03918_ _04092_ _04093_ _03866_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06264_ _01728_ _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05215_ _00769_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08003_ _01791_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10966__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06195_ _01359_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08577__A1 _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ delay_cycles\[14\] _04846_ _04843_ _04536_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08905_ _03959_ _03969_ _03982_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09885_ _04505_ _04792_ _04795_ net56 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10136__A1 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07001__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10270__I _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07065__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _03914_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05364__I _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08767_ _03758_ _03859_ _03865_ net147 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09829__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05979_ _01398_ _01522_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11018__D _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07718_ _02984_ _02991_ _02993_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08675__I _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ _03201_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08501__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ mem.mem_dff.code_mem\[30\]\[3\] _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10496__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06195__I _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10660_ _00252_ clknet_leaf_78_clock mem.mem_dff.code_mem\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__A2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09319_ _04266_ _04297_ _04300_ _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06115__I0 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10591_ _00183_ clknet_leaf_87_clock mem.mem_dff.code_mem\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08804__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06815__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08568__A1 _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _00735_ clknet_leaf_156_clock stack\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06043__A2 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11121__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11074_ _00666_ clknet_leaf_40_clock wb_write_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10127__A1 _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10025_ _04884_ _04896_ _04897_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10839__CLK clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08585__I _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09296__A2 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ _00519_ clknet_leaf_148_clock stack\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _00450_ clknet_leaf_168_clock stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10989__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10789_ _00381_ clknet_leaf_159_clock stack\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06806__A1 _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__C _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08253__C _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__A2 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09220__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10366__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__B _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05468__S1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _02391_ _02385_ _02392_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10118__A1 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10118__B2 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ _00777_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09670_ _04598_ _04629_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06882_ mem.mem_dff.code_mem\[9\]\[5\] _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08621_ _03744_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05833_ _01303_ _01375_ _01376_ _01298_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ _03705_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05764_ _01299_ _01300_ _01301_ _01304_ _01307_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_82_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07503_ _02824_ _02819_ _02810_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08495__B1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08483_ _01764_ _03632_ _03651_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05695_ _01235_ _01237_ _01238_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_165_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ mem.mem_dff.code_mem\[24\]\[3\] _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09039__A2 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0_clock clknet_3_7_0_clock clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07365_ _02365_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09104_ _04061_ _04114_ _04132_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08798__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06316_ _01855_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07296_ _02651_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09035_ _04059_ _04067_ _04080_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06247_ _01743_ _01781_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11144__CLK clknet_leaf_177_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input66_I i_wb_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10357__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06178_ _01625_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09211__A2 _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07222__A1 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__A2 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09937_ delay_cycles\[9\] _04835_ _04832_ _04836_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10372__A4 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05784__A1 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05308__B _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09868_ _04784_ _04786_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08722__A1 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output222_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08722__B2 stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08819_ stack\[7\]\[0\] _03916_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09799_ _03098_ _04728_ _04738_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05536__B2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06918__I _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _00304_ clknet_leaf_29_clock mem.mem_dff.data_mem\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05839__A2 _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10643_ _00235_ clknet_leaf_120_clock mem.mem_dff.code_mem\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ _00166_ clknet_leaf_89_clock mem.mem_dff.code_mem\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07461__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09202__A2 _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10511__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08961__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _00718_ clknet_leaf_158_clock stack\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11057_ _00649_ clknet_leaf_23_clock delay_cycles\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10661__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08713__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__S _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10008_ _04883_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06828__I _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09204__I _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11017__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05480_ _01029_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06563__I mem.mem_dff.code_mem\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07150_ _02537_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06101_ _01578_ _01590_ _01204_ _01244_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07081_ _02376_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07452__A1 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06032_ _01575_ _01232_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10339__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__B _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05766__A1 _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07983_ _01616_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06231__C _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09722_ _04659_ _04681_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06934_ _02282_ _02367_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _04564_ _04566_ _04568_ _04562_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_55_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06865_ _02229_ _02324_ _02315_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05518__A1 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08604_ _03208_ _03748_ _03749_ net144 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05816_ _00769_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09584_ delay_cycles\[11\] _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06796_ _02149_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06191__A1 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _03690_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05747_ _01290_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08466_ _03635_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05678_ net134 _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07417_ _02754_ _02746_ _02757_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06494__A2 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08397_ _03581_ _03582_ _03583_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07348_ _02350_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07279_ _02648_ _02650_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07994__A2 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output172_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _03743_ _03940_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05844__I2 stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09196__B2 stack\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10684__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08943__A1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05221__A3 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09499__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05780__I1 stack\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09959__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08863__I _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _00218_ clknet_leaf_104_clock mem.mem_dff.code_mem\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10557_ _00149_ clknet_leaf_91_clock mem.mem_dff.code_mem\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05445__B1 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _00080_ clknet_leaf_99_clock mem.mem_dff.code_mem\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05996__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__B2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05727__I _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08103__I _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05748__A1 _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05748__B2 _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11109_ _00701_ clknet_leaf_141_clock stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09362__C _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06650_ _02138_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06173__A1 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05601_ _01138_ _01148_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06581_ _02095_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A1 stack\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _03505_ _03510_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05532_ stack\[14\]\[6\] _01080_ _01076_ stack\[15\]\[6\] _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08773__I _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05359__S0 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ mem.mem_dff.data_mem\[2\]\[3\] _03044_ _03375_ mem.mem_dff.data_mem\[6\]\[3\]
+ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ _01013_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07389__I mem.mem_dff.code_mem\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06507__B _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07202_ _02589_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08182_ _03015_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05394_ _00944_ _00945_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_146_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09414__A2 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07133_ _02532_ _02536_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__B1 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05838__S _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__B1 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07064_ _02436_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput210 net252 rambus_wb_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput221 net221 rambus_wb_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09178__A1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput232 net253 rambus_wb_we_o vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_161_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06015_ _00931_ _01557_ _01558_ _00891_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05637__I _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ mem.mem_dff.data_mem\[7\]\[5\] _03179_ _03176_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _04661_ _04662_ _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06917_ net240 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input29_I i_wb_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07897_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08153__A2 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _04583_ _04584_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06848_ _02309_ _02306_ _02310_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06468__I _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05372__I _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _04524_ _04525_ _04526_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06779_ _02170_ net230 _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_169_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08518_ _03198_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09498_ _00805_ _04449_ _04463_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07664__A1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _01630_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08861__B1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_185_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__A1 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10411_ _00003_ clknet_leaf_162_clock stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06931__I _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10342_ _03847_ _03662_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09169__B2 stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10273_ _05053_ _05098_ _05099_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08916__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08392__A2 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09689__I _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09644__A2 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10609_ _00201_ clknet_leaf_92_clock mem.mem_dff.code_mem\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07407__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08604__B1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05269__I0 stack\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08080__A1 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08907__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07820_ _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08383__A2 _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10190__A2 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ _03016_ _03018_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05992__I1 stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06702_ _02194_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A2 _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06288__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ _02962_ _02959_ _02964_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09883__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09421_ net153 _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06633_ _02102_ _02140_ _02130_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07894__A1 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05744__I1 stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09352_ mem.io_data_out\[5\] _04320_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06564_ _02072_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08303_ mem.mem_dff.code_mem\[7\]\[5\] _03428_ _02443_ mem.mem_dff.code_mem\[13\]\[5\]
+ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05515_ stack\[13\]\[5\] stack\[12\]\[5\] _00927_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09283_ _01172_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06495_ _02026_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08843__B1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08234_ mem.mem_dff.code_mem\[25\]\[3\] _02789_ _02846_ mem.mem_dff.code_mem\[27\]\[3\]
+ _03426_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05446_ stack\[11\]\[4\] stack\[8\]\[4\] stack\[9\]\[4\] stack\[10\]\[4\] _00953_
+ _00954_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_176_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05752__S0 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08165_ mem.mem_dff.code_mem\[17\]\[1\] _03358_ _03359_ mem.mem_dff.code_mem\[21\]\[1\]
+ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_181_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05377_ _00927_ stack\[0\]\[3\] stack\[1\]\[3\] _00928_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ _02059_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07949__A2 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ _02292_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07047_ _02224_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08359__C1 mem.mem_dff.code_mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05367__I _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__I _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08998_ _03712_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07949_ _03009_ _03162_ _03169_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output135_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__A1 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__B2 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _00552_ clknet_leaf_142_clock stack\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06137__A1 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__A2 _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07885__A1 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _04574_ _04489_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10891_ _00483_ clknet_leaf_0_clock stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09087__B1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05360__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08062__A1 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08062__B2 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10183__I _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10325_ _05132_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05277__I _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10116__C _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05820__B1 _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10256_ _01933_ _04016_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07706__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10187_ _04998_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06376__A1 _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10172__A2 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06376__B2 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05974__I1 stack\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07441__B _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05300_ _00772_ _00852_ _00853_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06280_ _01719_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06300__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05231_ net137 _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07667__I _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08053__A1 mem.io_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__B1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09970_ _04807_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05257__I3 stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09882__I _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08921_ _03827_ _03993_ _03994_ _03675_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_1_0_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _01640_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_133_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10163__A2 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07803_ _02943_ _03058_ _03054_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08783_ _01181_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05995_ stack\[14\]\[5\] stack\[15\]\[5\] _00770_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05965__I1 stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _02121_ _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10895__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__A2 _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _02949_ _02942_ _02950_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ _04367_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06616_ _02124_ _02115_ _02125_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _02840_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09608__A2 cycles_per_ms\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__I _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09335_ net104 _04304_ _02618_ net98 _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06547_ _02070_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input96_I rambus_wb_dat_i[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ net256 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06478_ mem.mem_dff.cycles\[1\] _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08217_ _03402_ _03408_ _03409_ _03410_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xclkbuf_leaf_180_clock clknet_4_4_0_clock clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05429_ _00980_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_58_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09278__B _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ _04177_ _04196_ _04201_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08148_ _02346_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09792__A1 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08079_ net74 _03273_ _03274_ net125 _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10110_ net178 _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11090_ _00682_ clknet_leaf_15_clock net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10041_ _04910_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10943_ _00535_ clknet_leaf_142_clock stack\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_clock clknet_4_6_0_clock clknet_leaf_133_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10874_ _00466_ clknet_leaf_178_clock stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06530__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11050__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10618__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__I _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07086__A2 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_148_clock clknet_4_5_0_clock clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10090__A1 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08035__A1 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__B1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08035__B2 stack\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10768__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09783__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08586__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09783__B2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10308_ _05123_ _05124_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08338__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__B _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _01643_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05735__I _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08889__A3 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09550__A4 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05947__I1 stack\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ stack\[24\]\[0\] stack\[25\]\[0\] _00792_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ _02613_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06401_ _01073_ _01907_ _01840_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07381_ mem.mem_dff.code_mem\[23\]\[0\] _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09877__I _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09120_ _03635_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06332_ _01025_ _01869_ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_176_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09051_ _04088_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06285__B1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06824__A2 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06263_ _00917_ _01773_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07397__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08002_ _03212_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05214_ _00768_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06194_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09774__A1 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08577__A2 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06588__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10384__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _04840_ _04848_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05260__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ _03842_ _03971_ _03979_ stack\[10\]\[4\] _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09884_ _04791_ _04796_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05645__I _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_clock clknet_3_5_0_clock clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ stack\[7\]\[4\] _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08956__I _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08766_ stack\[11\]\[3\] _03862_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_211_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05978_ stack\[18\]\[5\] stack\[19\]\[5\] stack\[16\]\[5\] stack\[17\]\[5\] _00800_
+ _00890_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I i_la_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_clock clknet_4_11_0_clock clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ mem.mem_dff.data_mem\[0\]\[0\] _02992_ _02982_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11073__CLK clknet_opt_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08697_ _01182_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08501__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _02935_ _02929_ _02937_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06476__I _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06512__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05380__I _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_65_clock clknet_4_11_0_clock clknet_leaf_65_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07579_ _02883_ _02878_ _02884_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _04263_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _00182_ clknet_leaf_87_clock mem.mem_dff.code_mem\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06115__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__A1 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _04169_ _04234_ _04240_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10072__B2 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10910__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08280__A4 _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05874__I0 stack\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A2 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05756__S _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11142_ _00734_ clknet_leaf_138_clock stack\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05251__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11073_ _00665_ clknet_opt_3_0_clock net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput110 reset net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10024_ delay_counter\[3\] _04888_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05929__I1 stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08866__I _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10926_ _00518_ clknet_leaf_147_clock stack\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05290__I _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ _00449_ clknet_leaf_168_clock stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10788_ _00380_ clknet_leaf_3_clock stack\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10063__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10590__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09205__B1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09756__A1 edge_interrupts vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10366__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__A1 exec.out_of_order_exec vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06950_ _02358_ _02386_ _02378_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I i_la_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05901_ _01275_ _01440_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06881_ _02333_ _02334_ _02336_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08620_ _03223_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05832_ stack\[30\]\[7\] stack\[31\]\[7\] _01371_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07680__I _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08551_ _03167_ _03704_ _03699_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05763_ _01306_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07502_ _02040_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08495__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ _03650_ _03642_ _03648_ stack\[19\]\[1\] _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08495__B2 stack\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05694_ _01224_ _01206_ _01229_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _02769_ _02764_ _02770_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10933__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08247__A1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07364_ _02702_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09400__I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09103_ _04131_ _04116_ _04127_ stack\[24\]\[5\] _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06315_ _01720_ _01833_ _01853_ _01854_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09995__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08798__A2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ _02651_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04011_ _04069_ _04078_ stack\[9\]\[4\] _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06246_ _00918_ _01746_ _01783_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10357__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input59_I i_wb_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__A2 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ delay_cycles\[9\] _04560_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_154_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10109__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05375__I _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05784__A2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09867_ _04537_ _04785_ _04780_ net48 _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08722__A2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10463__CLK clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08818_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06733__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09798_ net257 _04730_ _04731_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_46_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ stack\[11\]\[0\] _03862_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A1 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10711_ _00303_ clknet_leaf_30_clock mem.mem_dff.data_mem\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10642_ _00234_ clknet_leaf_103_clock mem.mem_dff.code_mem\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08238__A1 mem.mem_dff.code_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10573_ _00165_ clknet_leaf_81_clock mem.mem_dff.code_mem\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05311__I2 stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09738__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07213__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05224__A1 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _00717_ clknet_leaf_158_clock stack\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__A1 _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05285__I _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09980__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11056_ _00648_ clknet_leaf_24_clock delay_cycles\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06024__I0 stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08713__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ delay_counter\[0\] _04880_ _04882_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10956__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08477__A1 _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10284__A1 stack\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10909_ _00501_ clknet_leaf_139_clock stack\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08229__A1 mem.mem_dff.code_mem\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08229__B2 mem.mem_dff.code_mem\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06100_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ mem.mem_dff.code_mem\[14\]\[7\] _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__A1 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06031_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10339__A2 _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07675__I _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08401__A1 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08401__B2 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ _01605_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06963__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05766__A2 stack\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06933_ _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09721_ _04660_ _04665_ _04680_ _04388_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__B1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06864_ _02322_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09652_ _04610_ _04611_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06715__A1 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05518__A2 _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05815_ _01333_ _01339_ _01358_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08603_ _03744_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09583_ _04488_ _04534_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06020__S _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06795_ mem.mem_dff.code_mem\[7\]\[3\] _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _01711_ _03674_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05746_ _01280_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ _03634_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05677_ _01200_ _01213_ _01220_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08455__B intr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07416_ _02755_ _02747_ _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ net121 _03107_ _03578_ _03579_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07347_ _02702_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07278_ _02649_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_opt_4_1_clock_I clknet_opt_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _03989_ _03824_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06229_ _01556_ _01571_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05844__I3 stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09196__A2 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09735__A4 cycles_per_ms\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08943__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05319__B _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _04805_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06006__I0 stack\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A3 _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_181_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09305__I _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10266__A1 _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07131__A1 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06664__I _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05693__A1 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10625_ _00217_ clknet_leaf_104_clock mem.mem_dff.code_mem\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10556_ _00148_ clknet_leaf_91_clock mem.mem_dff.code_mem\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08631__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05445__A1 stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05445__B2 _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10487_ _00079_ clknet_leaf_118_clock mem.mem_dff.code_mem\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05996__A2 _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11108_ _00700_ clknet_leaf_144_clock stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11039_ _00631_ clknet_leaf_33_clock cycles_per_ms\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07444__B _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06173__A2 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ _01127_ _01143_ _01147_ _01053_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06580_ _02020_ net229 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10257__A1 stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05531_ _01049_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05359__S1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08250_ mem.mem_dff.code_mem\[0\]\[3\] _03290_ _03434_ _03442_ _03316_ _03443_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_20_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06574__I mem.mem_dff.code_mem\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05462_ _00855_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07201_ _02532_ _02588_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08181_ mem.mem_dff.data_mem\[2\]\[1\] _03044_ _03375_ mem.mem_dff.data_mem\[6\]\[1\]
+ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10096__I _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05393_ _00801_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__A4 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07132_ _02535_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08622__B2 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05436__A1 stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ mem.mem_dff.code_mem\[14\]\[3\] _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05436__B2 stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput200 net200 rambus_wb_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput211 net248 rambus_wb_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput222 net222 rambus_wb_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06014_ stack\[2\]\[1\] stack\[3\]\[1\] _01463_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09178__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07965_ _03001_ _03178_ _03180_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09704_ _04663_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06749__I mem.mem_dff.code_mem\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06916_ _02348_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ _03131_ _03017_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05653__I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ _04588_ _04591_ _04594_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06847_ _02246_ _02307_ _02303_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07361__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09566_ _04522_ _04521_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06778_ mem.mem_dff.code_mem\[7\]\[0\] _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10501__CLK clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05729_ _00941_ stack\[7\]\[2\] _01272_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08517_ _03678_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07113__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09497_ _02000_ _04462_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08310__B1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08861__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ _03616_ _01696_ _03618_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08861__B2 stack\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05675__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08379_ _03567_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_128_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10410_ _00002_ clknet_leaf_139_clock stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10651__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05278__I1 stack\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10341_ _05064_ _05140_ _05147_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ _01793_ _05090_ _05095_ stack\[30\]\[1\] _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11007__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06659__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06155__A2 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08852__A1 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05666__A1 _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10608_ _00200_ clknet_leaf_92_clock mem.mem_dff.code_mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08604__A1 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08604__B2 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05269__I1 stack\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _00131_ clknet_leaf_98_clock mem.mem_dff.code_mem\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05738__I _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08907__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08383__A3 _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07750_ _03017_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05473__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06701_ _02128_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09332__A2 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _02963_ _02960_ _02953_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10524__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06632_ _02138_ _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09420_ _04386_ _04365_ _04393_ _04394_ _04375_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08784__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07894__A2 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06563_ mem.mem_dff.code_mem\[1\]\[4\] _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09351_ _04283_ mem.dff_data_out\[5\] _04330_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10966__D _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ mem.mem_dff.code_mem\[9\]\[5\] _03429_ _03432_ mem.mem_dff.code_mem\[14\]\[5\]
+ mem.mem_dff.code_mem\[28\]\[5\] _03430_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05514_ _00946_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10674__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09282_ _03241_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06494_ _02021_ _02025_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08843__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08843__B2 stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08233_ _03425_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05445_ stack\[14\]\[4\] _00925_ _00946_ _00995_ _00921_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_147_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05752__S1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05849__S _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08164_ _02675_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08225__S _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05376_ _00902_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ mem.mem_dff.code_mem\[15\]\[6\] _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ mem.mem_dff.code_mem\[23\]\[0\] _02731_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05648__I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07046_ mem.mem_dff.code_mem\[14\]\[0\] _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08959__I _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__A1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input41_I i_wb_addr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ _04050_ _04052_ _04053_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07582__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ mem.mem_dff.data_mem\[6\]\[7\] _03163_ _03168_ _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_54_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09323__A2 _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _03115_ _03116_ _03118_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output128_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09618_ _04572_ _04573_ _04576_ _04577_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07885__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10890_ _00482_ clknet_leaf_183_clock stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05896__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ delay_cycles\[16\] _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09087__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09087__B2 stack\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07103__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06860__A3 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10324_ stack\[16\]\[0\] _05135_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06073__A1 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05820__A1 _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10255_ _05064_ _05071_ _05085_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05820__B2 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09011__A1 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05259__S0 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10547__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _05031_ _05033_ _05034_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05293__I _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05584__B1 stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09314__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10697__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05887__A1 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09078__A1 stack\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05887__B2 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08825__A1 stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06300__A2 _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05230_ net135 _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09250__A1 _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__B2 stack\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06064__A1 _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08920_ _01690_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__I mem.mem_dff.code_mem\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08851_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07802_ _03045_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_5_0_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05994_ stack\[12\]\[5\] stack\[13\]\[5\] _01410_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08782_ _03887_ _03885_ _03871_ _03856_ _03888_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08108__A3 _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ _03001_ _03002_ _03004_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07316__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ _02867_ _02944_ _02939_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09403_ _04376_ _04378_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06615_ _02060_ _02118_ _02112_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07595_ mem.mem_dff.code_mem\[28\]\[7\] _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06546_ _02025_ _02069_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09334_ _04264_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08816__A1 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06477_ _02009_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09265_ _04249_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_194_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06762__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08216_ mem.mem_dff.code_mem\[7\]\[2\] _02258_ _02469_ mem.mem_dff.code_mem\[14\]\[2\]
+ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05428_ _00949_ _00958_ _00978_ _00979_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA_input89_I rambus_wb_dat_i[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09196_ _04129_ _04186_ _04200_ stack\[20\]\[4\] _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08147_ mem.mem_dff.code_mem\[25\]\[1\] _03340_ _03341_ mem.mem_dff.code_mem\[27\]\[1\]
+ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05359_ stack\[7\]\[2\] stack\[4\]\[2\] stack\[5\]\[2\] stack\[6\]\[2\] _00811_ _00891_
+ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_175_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06055__A1 _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08078_ _03263_ _03277_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ _02394_ _02446_ _02453_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ delay_counter\[6\] _04909_ _04881_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06358__A2 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05566__B1 stack\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08504__B1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ _00534_ clknet_leaf_146_clock stack\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07858__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10873_ _00465_ clknet_leaf_149_clock stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08807__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09480__A1 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10090__A2 _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08035__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__B2 stack\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05288__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09783__A2 _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08991__B1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10307_ _03221_ _05109_ _05115_ _04103_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07717__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10238_ _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10143__B _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08743__B1 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__A4 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10169_ _04288_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05557__B1 _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06400_ _01936_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07380_ _02725_ _02716_ _02728_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05580__I0 stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06331_ _01024_ _01728_ _01867_ _01868_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08274__A2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09050_ _04085_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06285__A1 stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06285__B2 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06262_ _01740_ _01776_ _01802_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_148_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05332__I0 stack\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05213_ net135 _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08001_ _03210_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_198_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10712__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__A1 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ _01249_ _01731_ _01735_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06037__A1 _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ delay_cycles\[13\] _04846_ _04843_ _04847_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08903_ _03957_ _03970_ _03981_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05260__A2 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06023__S _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09883_ cycles_per_ms\[20\] _04792_ _04795_ net55 _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _03915_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08765_ _03875_ _03876_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05977_ _01380_ _01517_ _01520_ _01436_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _02990_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06757__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03736_ _03816_ _03818_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07647_ _02936_ _02931_ _02923_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ _02824_ _02879_ _02871_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09317_ _04298_ _04299_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06529_ _02055_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A1 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 exec.memory_input\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ _04218_ _04236_ _04238_ stack\[22\]\[1\] _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06276__B2 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output195_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05874__I1 stack\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ _04185_ _04186_ _04187_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06028__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11141_ _00733_ clknet_leaf_138_clock stack\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05836__I _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05251__A2 _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11072_ _00664_ clknet_leaf_87_clock net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput100 rambus_wb_dat_i[2] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10023_ _04894_ _04895_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08725__B1 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05539__B1 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06751__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10189__I _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10925_ _00517_ clknet_leaf_34_clock wb_read_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05504__C _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05306__A3 _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _00448_ clknet_leaf_162_clock stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10735__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09453__A1 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10787_ _00379_ clknet_leaf_3_clock stack\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10063__A2 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_176_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09205__A1 _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09205__B2 stack\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06019__A1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05947__S _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__B _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09218__I _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09508__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08122__I _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06990__A2 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05900_ _01401_ _01441_ _01443_ _01272_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06880_ _02242_ _02335_ _02331_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05831_ stack\[28\]\[7\] stack\[29\]\[7\] _01374_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09381__C _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05762_ _01305_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08550_ _03703_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05481__I _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ mem.mem_dff.code_mem\[26\]\[2\] _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08481_ _03214_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05693_ _01188_ _01198_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08495__A2 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09888__I _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07432_ _02710_ _02765_ _02756_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05702__B1 _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07363_ mem.mem_dff.code_mem\[22\]\[4\] _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09102_ _01922_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06314_ _01191_ _01820_ _01754_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07294_ mem.mem_dff.code_mem\[20\]\[4\] _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_202_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09033_ _04056_ _04068_ _04079_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06245_ _01761_ _01784_ _01786_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06176_ _01679_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07357__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_clock clknet_opt_6_0_clock clknet_leaf_132_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05656__I _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05233__A2 _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09935_ _04823_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08032__I _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11040__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _04768_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07871__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_147_clock clknet_4_5_0_clock clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08817_ _03185_ _03913_ _03914_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ _01795_ _04732_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07930__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06487__I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08748_ _03861_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05792__I0 stack\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09132__B1 _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output208_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ _03669_ _03807_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_4_9_0_clock clknet_3_4_0_clock clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _00302_ clknet_leaf_36_clock mem.mem_dff.data_mem\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10293__A2 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10641_ _00233_ clknet_leaf_103_clock mem.mem_dff.code_mem\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08238__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A1 _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10045__A2 _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _00164_ clknet_leaf_81_clock mem.mem_dff.code_mem\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09738__A2 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07749__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05855__S0 _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11124_ _00716_ clknet_leaf_158_clock stack\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11055_ _00647_ clknet_leaf_24_clock delay_cycles\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09482__B _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__I mem.mem_dff.data_mem\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09371__B1 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10006_ _04881_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06024__I1 stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08477__A2 _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10908_ _00500_ clknet_leaf_186_clock stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10284__A2 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10839_ _00431_ clknet_leaf_153_clock stack\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07988__A1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05838__I1 stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06030_ _01322_ _01573_ _01236_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06660__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05476__I _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07981_ _03186_ _03188_ _03189_ _03192_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_clock clknet_4_11_0_clock clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09720_ _04673_ _04675_ _04676_ _04679_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06932_ _02376_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07691__I mem.mem_dff.code_mem\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08165__B2 mem.mem_dff.code_mem\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__B1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09651_ _04544_ _04567_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06863_ _02322_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08602_ _03742_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05814_ _01279_ _01345_ _01350_ _01356_ _01357_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09582_ cycles_per_ms\[13\] _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05774__I0 stack\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06794_ _02266_ _02260_ _02267_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_clock clknet_4_15_0_clock clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08533_ _01893_ _03670_ _03689_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06100__I _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05745_ stack\[14\]\[2\] stack\[15\]\[2\] _00900_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07640__B _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input106_I rambus_wb_dat_i[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10275__A2 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08464_ _01673_ _01651_ _01679_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05676_ _01214_ _01215_ _01219_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09411__I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07415_ _02726_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__A1 _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ net121 _03573_ _03576_ _03107_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07346_ _02648_ _02701_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _02171_ _02534_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clock clknet_4_8_0_clock clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input71_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09016_ _03889_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06770__I mem.mem_dff.code_mem\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06228_ _01729_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06159_ _01700_ _01670_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10430__CLK clknet_leaf_75_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05386__I _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06403__A1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output158_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09918_ _04816_ _04822_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08697__I _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08156__A1 mem.mem_dff.code_mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_124_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__I1 stack\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _04354_ _04766_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10580__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06706__A2 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05765__I0 stack\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06945__I mem.mem_dff.code_mem\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A2 _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07131__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__I _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06166__B _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10624_ _00216_ clknet_leaf_104_clock mem.mem_dff.code_mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06890__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10555_ _00147_ clknet_leaf_95_clock mem.mem_dff.code_mem\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08631__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05445__A2 _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10486_ _00078_ clknet_leaf_119_clock mem.mem_dff.code_mem\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05296__I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__A1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08395__B2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10923__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11107_ _00699_ clknet_leaf_8_clock prev_reg_write vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08147__A1 mem.mem_dff.code_mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11038_ _00630_ clknet_leaf_33_clock cycles_per_ms\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06121__S _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09895__A1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05756__I0 stack\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10257__A2 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05530_ _01077_ stack\[12\]\[6\] stack\[13\]\[6\] _01078_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09231__I _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05461_ _01011_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ _02587_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ _03328_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05392_ _00883_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_220_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07131_ _02021_ _02534_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10453__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07686__I mem.mem_dff.code_mem\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06633__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06590__I mem.mem_dff.code_mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07062_ _02477_ _02471_ _02479_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05436__A2 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput201 net201 rambus_wb_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput212 net246 rambus_wb_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06013_ stack\[0\]\[1\] stack\[1\]\[1\] _01442_ _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput223 net223 rambus_wb_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_161_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10193__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07964_ mem.mem_dff.data_mem\[7\]\[4\] _03179_ _03176_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05995__I0 stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__B1 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09703_ _01800_ _01833_ _01959_ _04444_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06915_ mem.mem_dff.code_mem\[10\]\[4\] _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07895_ _03130_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09886__A1 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09634_ _04592_ _04580_ _04582_ _04593_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06846_ mem.mem_dff.code_mem\[8\]\[5\] _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09565_ delay_cycles\[19\] _04510_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06777_ _02250_ _02241_ _02253_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10248__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _01707_ _03200_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_212_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05728_ _01271_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _04440_ _01615_ _04451_ _04461_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08310__A1 mem.mem_dff.code_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08447_ _01664_ _03617_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05659_ _01198_ _01200_ _01202_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08861__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__I _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ mem.dff_data_out\[7\] _03566_ _03483_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07329_ _02677_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__A1 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08613__A2 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07596__I _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05278__I2 stack\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _01923_ _05132_ _05145_ stack\[16\]\[5\] _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10946__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _05097_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08377__A1 _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__A1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__I _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05780__S _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06675__I _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08301__A1 mem.mem_dff.code_mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_6_0_clock clknet_2_3_0_clock clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10476__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__I _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__I _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _00199_ clknet_leaf_92_clock mem.mem_dff.code_mem\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08604__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06615__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _00130_ clknet_leaf_113_clock mem.mem_dff.code_mem\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10146__B _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10469_ _00061_ clknet_leaf_56_clock mem.mem_dff.code_mem\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08368__A1 _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07040__A1 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08383__A4 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11101__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09868__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ mem.mem_dff.code_mem\[4\]\[7\] _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ _02036_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08540__A1 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06631_ _02138_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05354__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09350_ _04328_ _04329_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06562_ _02080_ _02073_ _02082_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10819__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08301_ mem.mem_dff.code_mem\[25\]\[5\] _02789_ _02846_ mem.mem_dff.code_mem\[27\]\[5\]
+ _03491_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05513_ stack\[15\]\[5\] _01062_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09281_ _03622_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06493_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08843__A2 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ mem.mem_dff.code_mem\[10\]\[3\] _02347_ _02762_ mem.mem_dff.code_mem\[24\]\[3\]
+ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05444_ stack\[13\]\[4\] stack\[12\]\[4\] _00942_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__CLK clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08163_ _02561_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05375_ _00926_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _02519_ _02516_ _02520_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08094_ _03289_ _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02463_ _02456_ _02465_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08359__A1 mem.mem_dff.code_mem\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10166__A1 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _04004_ _04048_ _04046_ stack\[25\]\[1\] _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I i_wb_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _03167_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09859__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__B2 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ _03086_ _03117_ _03113_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09617_ cycles_per_ms\[6\] _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06829_ _02229_ _02296_ _02283_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05345__A1 _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10499__CLK clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09548_ _04485_ _04495_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05896__A2 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08295__B1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _04403_ _03199_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08598__A1 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10323_ _05134_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06073__A2 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11124__CLK clknet_leaf_158_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10254_ _04227_ _05073_ _05082_ stack\[14\]\[5\] _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05820__A2 _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09011__A2 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07022__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05259__S1 _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10185_ _04288_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05959__I0 stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05574__I _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__A2 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05584__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05584__B2 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A1 _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09078__A2 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08825__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08125__I _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09250__A2 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07261__A1 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10148__A1 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07013__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10390__I _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08210__B1 _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08850_ _03939_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07801_ _03045_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08761__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ stack\[11\]\[7\] _03872_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05993_ _01426_ _01535_ _01536_ _01430_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07732_ mem.mem_dff.data_mem\[0\]\[4\] _03003_ _02999_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10641__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07663_ mem.mem_dff.code_mem\[30\]\[6\] _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10320__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09402_ exec.out_of_order_exec _04359_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06614_ mem.mem_dff.code_mem\[2\]\[6\] _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07594_ _02894_ _02889_ _02895_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09069__A2 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09333_ _01227_ _04265_ _04314_ _04289_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06545_ _02019_ net228 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10791__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08816__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09264_ net143 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06476_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08215_ mem.mem_dff.code_mem\[9\]\[2\] _02321_ _02876_ mem.mem_dff.code_mem\[28\]\[2\]
+ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05427_ _00854_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09195_ _04188_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_194_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08146_ _02845_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05358_ _00910_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10387__A1 _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06055__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ mem.io_data_out\[4\] _03267_ _03271_ _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05289_ _00810_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07028_ _02436_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__C _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07004__A1 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output140_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05566__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _01932_ _03235_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05566__B2 _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07823__B _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__A1 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08504__B2 stack\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10941_ _00533_ clknet_leaf_0_clock stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10311__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05343__B _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _00464_ clknet_leaf_152_clock stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08807__A2 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06953__I _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09469__C _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09232__A2 _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10514__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07784__I _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10306_ stack\[27\]\[3\] _05112_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08991__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__B2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05518__B _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10237_ _03635_ _03701_ _03994_ _03945_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_79_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08743__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__B2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _04540_ _05020_ _05013_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05557__A1 stack\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05557__B2 stack\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10099_ _00877_ _04928_ _04965_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09504__I _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10302__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05580__I1 stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07959__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06330_ _01867_ _01868_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06863__I _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_2_3_0_clock clknet_0_clock clknet_2_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07482__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__A2 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10385__I stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ _01782_ _01775_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05332__I1 stack\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05479__I _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08000_ _03206_ _03211_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_204_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05212_ _00766_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10369__A1 _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06192_ _01732_ _01634_ _01734_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09223__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_97_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07785__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08982__A1 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ delay_cycles\[13\] _04534_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08902_ _03839_ _03972_ _03979_ stack\[10\]\[3\] _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09882_ _04774_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A1 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08833_ _03926_ _03927_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05548__A1 stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__C _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05399__I1 stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07643__B _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _03755_ _03864_ _03865_ net146 _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05976_ _01467_ _01518_ _01519_ _01298_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07715_ _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ _03696_ _03801_ _03813_ stack\[5\]\[7\] _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _02040_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ mem.mem_dff.code_mem\[28\]\[2\] _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _01800_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06528_ net237 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09462__A2 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10537__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _04066_ _04234_ _04239_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06459_ _00763_ _01172_ _01993_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_182_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05389__I _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _03202_ _04086_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output188_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _02290_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06028__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__B _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10687__CLK clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11140_ _00732_ clknet_leaf_138_clock stack\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_clock clknet_3_2_0_clock clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_122_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11071_ _00663_ clknet_opt_5_0_clock net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput101 rambus_wb_dat_i[30] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08725__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10022_ delay_counter\[3\] _04649_ _04885_ _00983_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05539__A1 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05539__B2 stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__B1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ _00516_ clknet_leaf_186_clock stack\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _00447_ clknet_leaf_160_clock stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10786_ _00378_ clknet_leaf_170_clock stack\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07464__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10063__A3 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_119_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09205__A2 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07216__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10154__B _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05963__S _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05830_ _00820_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06858__I _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05761_ _00773_ _01270_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ _02821_ _02817_ _02822_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10287__B1 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _01183_ _03632_ _03649_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05692_ _01193_ _01234_ _01219_ _01235_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07431_ mem.mem_dff.code_mem\[24\]\[2\] _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ _02712_ _02703_ _02714_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _04059_ _04114_ _04130_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06313_ _01801_ _01845_ _01849_ _01852_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06258__A2 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07293_ _02659_ _02652_ _02661_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05305__I1 stack\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08652__B1 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ _04008_ _04070_ _04078_ stack\[9\]\[3\] _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06244_ _00876_ _01785_ _01782_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06175_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_172_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06542__B _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05313__S0 _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ _04829_ _04834_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06430__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08707__A1 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09865_ _03281_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _03645_ _03807_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09796_ _00756_ _04728_ _04736_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05672__I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07930__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _03740_ _03859_ _03860_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05959_ stack\[2\]\[4\] stack\[3\]\[4\] stack\[0\]\[4\] stack\[1\]\[4\] _00868_ _00869_
+ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05605__C _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09132__B2 stack\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08678_ _03772_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__C1 mem.mem_dff.code_mem\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07629_ mem.mem_dff.code_mem\[29\]\[7\] _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07694__A1 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _00232_ clknet_leaf_103_clock mem.mem_dff.code_mem\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06249__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _00163_ clknet_leaf_81_clock mem.mem_dff.code_mem\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_120_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__C _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09738__A3 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07749__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08946__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05304__S0 _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11123_ _00715_ clknet_leaf_192_clock stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06421__A2 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05855__S1 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08961__A4 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11054_ _00646_ clknet_leaf_25_clock delay_cycles\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09371__A1 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10005_ _04640_ _04645_ _04805_ _01644_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09371__B2 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07921__A2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A3 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _00499_ clknet_leaf_186_clock stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10838_ _00430_ clknet_leaf_154_clock stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10852__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06119__S _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07302__I mem.mem_dff.code_mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__B _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10769_ _00361_ clknet_leaf_31_clock net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07980_ _03190_ _03191_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06931_ _02127_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09362__B2 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ cycles_per_ms\[11\] _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06862_ _02286_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clock clock clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05492__I _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ stack\[3\]\[0\] _03746_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05813_ _00777_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09581_ _04486_ _04530_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06793_ _02235_ _02261_ _02252_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05774__I1 stack\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _03659_ _03676_ _03687_ stack\[29\]\[5\] _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05744_ stack\[12\]\[2\] stack\[13\]\[2\] _00857_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__A3 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08463_ _01757_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10985__D _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05675_ _01216_ _01218_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07414_ _02526_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08394_ _03568_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08625__B1 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ _02531_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09015_ _04019_ _04063_ _04051_ _03987_ _04065_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_152_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06227_ net54 _01765_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_163_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08928__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input64_I i_wb_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06158_ _01700_ _01619_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06089_ _01632_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09917_ _04574_ _04811_ _04820_ _04821_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10725__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05616__B _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09848_ _04356_ _04759_ _04773_ _03569_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output220_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09779_ _04468_ _01179_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05765__I1 stack\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10875__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__B1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07122__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10623_ _00215_ clknet_leaf_104_clock mem.mem_dff.code_mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08616__B1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05778__S _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10554_ _00146_ clknet_leaf_80_clock mem.mem_dff.code_mem\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08092__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10485_ _00077_ clknet_leaf_56_clock mem.mem_dff.code_mem\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05577__I _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09592__A1 _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09493__B _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__I _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_2_0_clock clknet_2_1_0_clock clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_2_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_193_clock clknet_4_1_0_clock clknet_leaf_193_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11106_ _00698_ clknet_leaf_35_clock net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11037_ _00629_ clknet_leaf_33_clock cycles_per_ms\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06158__A1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__A2 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout251_I net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_131_clock clknet_4_6_0_clock clknet_leaf_131_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08128__I _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05460_ _01010_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05391_ stack\[5\]\[3\] stack\[4\]\[3\] _00942_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_clock clknet_4_5_0_clock clknet_leaf_146_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_199_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07061_ _02478_ _02473_ _02464_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07830__A1 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput202 net202 rambus_wb_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06012_ _01548_ _01555_ _01424_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput213 net243 rambus_wb_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput224 net224 rambus_wb_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09032__B1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__A2 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05444__I0 stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07963_ _03170_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05995__I1 stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__A1 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09335__B2 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06914_ _02360_ _02349_ _02362_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09702_ _01800_ _01833_ _01960_ _04444_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07894_ _02020_ _03014_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06845_ _02305_ _02306_ _02308_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09633_ cycles_per_ms\[4\] _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06111__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07651__B _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09564_ cycles_per_ms\[19\] _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06776_ _02165_ _02243_ _02252_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _03676_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05727_ _01270_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09495_ _04441_ _01613_ _04460_ _04339_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_169_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08310__A2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _01662_ _01663_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05658_ _01201_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08377_ _03560_ _03565_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05589_ _01089_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07328_ mem.mem_dff.code_mem\[21\]\[4\] _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _02621_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05278__I3 stack\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _05093_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output170_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__B _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06730__B _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__A2 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08376__C _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11053__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__B1 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__B2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06691__I _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10606_ _00198_ clknet_leaf_92_clock mem.mem_dff.code_mem\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08065__A1 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09262__B1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10537_ _00129_ clknet_leaf_113_clock mem.mem_dff.code_mem\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05823__B1 _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_78_clock clknet_4_15_0_clock clknet_leaf_78_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10468_ _00060_ clknet_leaf_56_clock mem.mem_dff.code_mem\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10399_ _03724_ _05172_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08411__I _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__B _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05971__S _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06630_ _02018_ _02137_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08540__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_clock clknet_4_2_0_clock clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06551__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05354__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05985__S0 _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06561_ _02045_ _02074_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08300_ _03490_ _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05512_ _00993_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10420__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09280_ _04264_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06492_ _02022_ _02023_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06303__A1 _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08231_ mem.mem_dff.code_mem\[8\]\[3\] _02293_ _02701_ mem.mem_dff.code_mem\[22\]\[3\]
+ _03423_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_220_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05443_ stack\[15\]\[4\] _00993_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06815__B _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ mem.mem_dff.code_mem\[1\]\[1\] _03355_ _02535_ mem.mem_dff.code_mem\[16\]\[1\]
+ _03356_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_159_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08056__A1 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09253__B1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05374_ _00881_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_167_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10570__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _02489_ _02517_ _02513_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07803__A1 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ _02290_ _02987_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05814__B1 _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ _02407_ _02457_ _02464_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08359__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10166__A2 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08995_ _04051_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ _01998_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06790__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__A2 _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I i_wb_addr[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ _03102_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A2 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09616_ delay_cycles\[6\] _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06828_ _02294_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06542__A1 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06759_ _02237_ _02228_ _02239_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09547_ cycles_per_ms\[18\] _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09478_ _04440_ _04446_ _04439_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08429_ net114 _03603_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10913__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09795__A1 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08598__A2 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _05075_ _05132_ _05133_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06073__A3 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__C _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10253_ _05061_ _05071_ _05084_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07022__A2 _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _04524_ _05032_ _05025_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05959__I1 stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06781__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05584__A2 stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09490__C _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08387__B _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08522__A2 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06686__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08286__B2 mem.mem_dff.data_mem\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10593__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__A1 single_step vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__I0 stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__B1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05966__S _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07013__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07800_ mem.mem_dff.data_mem\[2\]\[4\] _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08761__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08780_ _03853_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05992_ stack\[8\]\[5\] stack\[9\]\[5\] _01427_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07731_ _02990_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09710__A1 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _02946_ _02942_ _02948_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_93_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06613_ _02120_ _02115_ _02123_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04376_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _02867_ _02890_ _02886_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10936__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06544_ mem.mem_dff.code_mem\[1\]\[0\] _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09332_ _04303_ _04311_ _04313_ _04301_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10084__A1 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09263_ _04205_ _04246_ _04248_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_205_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06475_ _01997_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_205_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _03403_ _03404_ _03406_ _03407_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05426_ _00967_ _00971_ _00975_ _00977_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09226__B1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09194_ _04175_ _04196_ _04199_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07220__I _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__I2 stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _02788_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09777__A1 single_step vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05357_ stack\[3\]\[2\] stack\[0\]\[2\] stack\[1\]\[2\] stack\[2\]\[2\] _00901_ _00902_
+ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10387__A2 _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ net116 _03272_ _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05288_ _00842_ net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07027_ mem.mem_dff.code_mem\[13\]\[3\] _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08201__A1 mem.mem_dff.code_mem\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05608__C _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10466__CLK clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05566__A2 stack\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08978_ _03731_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07929_ mem.mem_dff.data_mem\[6\]\[0\] _03156_ _03152_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output133_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09701__A1 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10940_ _00532_ clknet_leaf_191_clock stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05318__A2 _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10311__A2 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10871_ _00463_ clknet_leaf_145_clock stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_1_0_clock clknet_3_0_0_clock clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08440__A1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09485__C _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10305_ _05121_ _05122_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08991__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05585__I _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10809__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10236_ _05071_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10167_ _04976_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06754__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05557__A2 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10098_ _04959_ _04960_ _04962_ _04964_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10959__CLK clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_1_0_clock_I clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10302__A2 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07305__I mem.mem_dff.code_mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05580__I2 stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06260_ _01729_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05332__I2 stack\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05211_ net136 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06191_ _01225_ _01733_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07975__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08431__A1 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09950_ _04823_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06993__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05495__I _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _03954_ _03970_ _03980_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _04791_ _04794_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _03758_ _03913_ _03920_ net147 _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__B _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05548__A2 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05399__I2 stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08763_ stack\[11\]\[2\] _03862_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05975_ stack\[30\]\[5\] stack\[31\]\[5\] _01371_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_211_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07714_ _02985_ _02986_ _02989_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08694_ _03732_ _03816_ _03817_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07215__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ mem.mem_dff.code_mem\[30\]\[2\] _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07170__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11114__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07576_ _02881_ _02878_ _02882_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__I _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10057__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06527_ mem.mem_dff.code_mem\[0\]\[5\] _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09315_ _03621_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09998__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input94_I rambus_wb_dat_i[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08046__I _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06458_ _01177_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09246_ _01758_ _04236_ _04238_ stack\[22\]\[0\] _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_210_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05484__A1 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05409_ _00887_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05484__B2 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ _04145_ _04025_ _03777_ _03233_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06389_ _01677_ _01925_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _03130_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08059_ _02002_ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11070_ _00662_ clknet_leaf_69_clock net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10021_ _04890_ _04891_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput102 rambus_wb_dat_i[31] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08725__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07834__B _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05539__A2 stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08489__A1 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__B2 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10923_ _00515_ clknet_leaf_187_clock stack\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10854_ _00446_ clknet_leaf_160_clock stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10048__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10785_ _00377_ clknet_leaf_169_clock stack\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_41_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10631__CLK clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08413__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__A1 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10781__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _04222_ _05050_ _05048_ stack\[12\]\[3\] _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11199_ net233 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06727__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10170__B _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05760_ _01303_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10287__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05691_ net130 net129 _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ _02767_ _02764_ _02768_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06874__I _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05702__A2 _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07361_ _02631_ _02705_ _02713_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10396__I _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08247__A4 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09100_ _04129_ _04116_ _04127_ stack\[24\]\[4\] _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06312_ _01814_ _01808_ _01850_ _01835_ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_07292_ _02631_ _02653_ _02660_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__A1 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05305__I2 stack\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08652__B2 stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09031_ _04073_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05466__A1 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06243_ _01226_ _01749_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06174_ _01644_ _01714_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08955__A2 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05313__S1 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09933_ _04555_ _04824_ _04832_ _04833_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08707__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09864_ _04783_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06718__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09425__I _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09380__A2 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ _03741_ _03637_ _01930_ _03640_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ _04376_ _04730_ _04731_ _04735_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07391__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08746_ _03743_ _03823_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05958_ _01485_ stack\[6\]\[4\] _01434_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10278__A1 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__A2 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05889_ stack\[14\]\[6\] stack\[15\]\[6\] _00827_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ _03804_ _03806_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__B1 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08340__C2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _02920_ _02915_ _02921_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07559_ _02866_ _02861_ _02868_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10654__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10570_ _00162_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05457__A1 _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09229_ _04225_ _04210_ _04223_ stack\[21\]\[4\] _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06733__B _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09738__A4 _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05209__A1 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10202__A1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A2 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05304__S1 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11122_ _00714_ clknet_leaf_189_clock stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06009__I0 stack\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11053_ _00645_ clknet_leaf_25_clock delay_cycles\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06709__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10004_ delay_counter\[0\] _04647_ _04879_ _00841_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09371__A2 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A2 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__B1 _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10906_ _00498_ clknet_leaf_185_clock stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__A1 stack\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05240__S0 _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _00429_ clknet_leaf_139_clock stack\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08634__A1 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ _00360_ clknet_leaf_31_clock net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _00291_ clknet_leaf_66_clock mem.mem_dff.data_mem\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__B _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05974__S _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06930_ mem.mem_dff.code_mem\[10\]\[7\] _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I i_la_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08289__C _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__A2 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06861_ _02320_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10527__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _03745_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05812_ _01267_ _01351_ _01354_ _01342_ _01355_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_95_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09580_ cycles_per_ms\[15\] _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06792_ mem.mem_dff.code_mem\[7\]\[2\] _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05743_ _01011_ _01283_ _01284_ _01286_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08531_ _01861_ _03670_ _03688_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08462_ _03631_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05674_ _01217_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05687__A1 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ mem.mem_dff.code_mem\[23\]\[7\] _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08393_ _03569_ _03577_ _03580_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05441__C _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07344_ _02467_ _02534_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08625__A1 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09848__C _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08625__B2 stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05439__A1 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05439__B2 stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07275_ mem.mem_dff.code_mem\[20\]\[0\] _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09014_ stack\[25\]\[7\] _04046_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08640__A4 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06226_ _01766_ _01767_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08928__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _01113_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05884__S _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input57_I i_wb_data[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _01622_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09916_ _04582_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05611__B2 stack\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09889__B1 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09155__I _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _04572_ _04757_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _03623_ _04475_ _04722_ _04708_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_46_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _03794_ _03825_ _03845_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06728__B _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10030__S _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__B2 stack\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07403__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05517__I2 stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11072__D _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10622_ _00214_ clknet_leaf_104_clock mem.mem_dff.code_mem\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08616__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08616__B2 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10553_ _00145_ clknet_leaf_80_clock mem.mem_dff.code_mem\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10484_ _00076_ clknet_leaf_56_clock mem.mem_dff.code_mem\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09041__A1 stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__C _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _00697_ clknet_leaf_35_clock net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05593__I _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11036_ _00628_ clknet_leaf_32_clock cycles_per_ms\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06158__A2 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05669__A1 _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05390_ _00941_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_159_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07060_ _02357_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06011_ _01408_ _01551_ _01554_ _01422_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_127_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput203 net203 rambus_wb_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09032__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput214 net240 rambus_wb_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09032__B2 stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput225 net225 rambus_wb_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07983__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05444__I1 stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06599__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07962_ _03170_ _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ _01769_ _04325_ _01896_ _01988_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09335__A2 _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06913_ _02269_ _02352_ _02361_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07346__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07893_ mem.mem_dff.data_mem\[5\]\[0\] _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09632_ cycles_per_ms\[5\] _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_163_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06844_ _02242_ _02307_ _02303_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09563_ _04519_ _04520_ _04521_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06775_ _02251_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08514_ _03672_ _03673_ _03189_ _03675_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_05726_ net137 _00775_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_64_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ _04442_ _04312_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08445_ _01660_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05657_ _01184_ _01185_ _01187_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08376_ mem.mem_dff.data_mem\[0\]\[7\] _03475_ _03476_ _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05588_ _01129_ _01132_ _01135_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10405__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07327_ _02685_ _02678_ _02687_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05678__I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A1 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ mem.mem_dff.code_mem\[19\]\[4\] _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06209_ _01225_ _01748_ _01750_ _01751_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07189_ _02578_ _02575_ _02579_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09023__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output163_I net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__B1 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06302__I _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__A1 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11067__D _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10992__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__B2 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06312__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10605_ _00197_ clknet_leaf_93_clock mem.mem_dff.code_mem\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09262__A1 _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09262__B2 stack\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06076__A1 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10536_ _00128_ clknet_leaf_115_clock mem.mem_dff.code_mem\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05823__A1 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 stack\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05823__B2 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10467_ _00059_ clknet_leaf_57_clock mem.mem_dff.code_mem\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08368__A3 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10398_ _05186_ _05170_ _05187_ _05189_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06379__A2 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05587__B1 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ _00611_ clknet_leaf_7_clock cycles_per_ms\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07879__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06000__A1 _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05985__S1 _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ _02065_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08828__A1 stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05511_ _01057_ _01058_ _01060_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06491_ net254 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08230_ _03420_ _03421_ _03422_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05442_ _00959_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10715__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _02026_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05373_ _00924_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09253__B2 stack\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07112_ mem.mem_dff.code_mem\[15\]\[5\] _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ _03282_ _03288_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07043_ _02436_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05814__A1 _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__I _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__A1 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__B1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05447__B _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08994_ _03669_ _03941_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__C _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07945_ _03007_ _03162_ _03166_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07319__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ _03102_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09433__I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09615_ delay_cycles\[5\] _04574_ _04489_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06827_ _02294_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _04500_ _04501_ _04504_ _04505_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06758_ _02150_ _02230_ _02238_ _02239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08819__A1 stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05709_ _01236_ _01240_ _01252_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09477_ _01700_ _04441_ _04445_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06689_ mem.mem_dff.code_mem\[4\]\[4\] _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07888__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08428_ _02037_ _03602_ _03606_ _03605_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_192_clock clknet_4_1_0_clock clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05353__I0 stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08047__A2 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ mem.mem_dff.code_mem\[7\]\[7\] _02257_ _03429_ mem.mem_dff.code_mem\[9\]\[7\]
+ mem.mem_dff.code_mem\[28\]\[7\] _02875_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05805__A1 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _03202_ _03643_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05281__A2 _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10252_ _04225_ _05073_ _05082_ stack\[14\]\[4\] _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07558__A1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _04976_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05959__I2 stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11020__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06781__A2 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07572__B _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_1_0_clock_I clknet_2_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_145_clock clknet_4_5_0_clock clknet_leaf_145_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09483__A1 _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06297__A1 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10093__A2 _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__A1 _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05895__I1 stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__B2 stack\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06049__A1 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10888__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10519_ _00111_ clknet_leaf_112_clock mem.mem_dff.code_mem\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08422__I _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07013__A3 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05991_ stack\[10\]\[5\] stack\[11\]\[5\] _01463_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08349__I0 mem.dff_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06772__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ _02990_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ _02947_ _02944_ _02939_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09710__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07721__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ net139 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06612_ _02122_ _02118_ _02112_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07592_ mem.mem_dff.code_mem\[28\]\[6\] _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ _04298_ _04312_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06543_ _02062_ _02049_ _02067_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__A2 _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ _04206_ _04232_ _04242_ stack\[22\]\[7\] _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05335__I0 _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06474_ _02005_ _02007_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08213_ mem.mem_dff.code_mem\[17\]\[2\] _03358_ _02620_ mem.mem_dff.code_mem\[19\]\[2\]
+ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05425_ _00922_ _00976_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ _04126_ _04192_ _04189_ stack\[20\]\[3\] _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09226__B2 stack\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__I3 stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ mem.mem_dff.code_mem\[7\]\[1\] _02258_ _02469_ mem.mem_dff.code_mem\[14\]\[1\]
+ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09777__A2 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05356_ _00889_ _00904_ _00907_ _00908_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09856__C _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07788__A1 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07657__B _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08075_ net73 _03273_ _03274_ net124 _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05287_ _00841_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07026_ _02450_ _02445_ _02451_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06212__A1 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _03961_ _04022_ _04037_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_62_clock clknet_4_14_0_clock clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07960__A1 mem.mem_dff.data_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07928_ _03154_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09162__B1 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output126_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ _03102_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A1 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10102__I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10870_ _00462_ clknet_leaf_152_clock stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_77_clock clknet_4_14_0_clock clknet_leaf_77_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ delay_cycles\[3\] delay_cycles\[2\] delay_cycles\[1\] delay_cycles\[0\] _04489_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08268__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__B1 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_clock clknet_4_8_0_clock clknet_leaf_15_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_193_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10304_ _03218_ _05114_ _05115_ _04100_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06451__A1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08728__B1 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10235_ _01640_ _03991_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10410__CLK clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ net167 _05011_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10097_ _04600_ _04963_ _04946_ intr\[1\] _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10560__CLK clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08900__B1 _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_5_0_clock_I clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10999_ _00591_ clknet_leaf_129_clock exec.memory_input\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05580__I3 stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10066__A2 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07321__I mem.mem_dff.code_mem\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05210_ _00765_ net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06190_ _01202_ _01245_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_204_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__B1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06442__A1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06993__A2 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ _03837_ _03972_ _03979_ stack\[10\]\[2\] _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09880_ _04524_ _04792_ _04788_ net53 _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ stack\[7\]\[3\] _03916_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10903__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05399__I3 stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08762_ _03869_ _03871_ _03873_ _03874_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05974_ stack\[28\]\[5\] stack\[29\]\[5\] _01438_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ _02014_ _02988_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08693_ _03694_ _03801_ _03813_ stack\[5\]\[6\] _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _02933_ _02929_ _02934_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07940__B _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ _02852_ _02879_ _02871_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09447__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _04267_ _04295_ _04296_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06526_ _02048_ _02049_ _02053_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10057__A2 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09245_ _04237_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06457_ _01934_ _01991_ _01992_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input87_I rambus_wb_dat_i[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05484__A2 stack\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05408_ _00959_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09176_ _03780_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06388_ _01684_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08127_ _03100_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05339_ stack\[19\]\[2\] stack\[16\]\[2\] stack\[17\]\[2\] stack\[18\]\[2\] _00843_
+ _00891_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10433__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09158__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06433__A1 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ _02005_ _03260_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06984__A2 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07009_ _02407_ _02429_ _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10020_ _04884_ _04892_ _04893_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput103 rambus_wb_dat_i[3] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10583__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07406__I mem.mem_dff.code_mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08489__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10296__A2 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10922_ _00514_ clknet_leaf_185_clock stack\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10853_ _00445_ clknet_leaf_160_clock stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06466__B _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10048__A2 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _00376_ clknet_leaf_159_clock stack\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A1 mem.mem_dff.code_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08110__B2 mem.mem_dff.code_mem\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05797__S _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06672__A1 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__A2 _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__A1 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05227__A2 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06424__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10220__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10926__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08177__A1 _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10218_ _03716_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11198_ net236 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07924__A1 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _05005_ _05006_ _04472_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06220__I _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07760__B _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10287__A2 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05690_ _01233_ _01215_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_208_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07360_ _02671_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06311_ _00982_ _01811_ _01835_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07291_ _02614_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__A2 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10456__CLK clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05305__I3 stack\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ _04054_ _04068_ _04077_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06242_ _01226_ _01634_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ _01618_ _01715_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06415__A1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04555_ _04557_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__A1 mem.mem_dff.code_mem\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08168__B2 mem.mem_dff.code_mem\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _04542_ _04769_ _04775_ net47 _03262_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08707__A3 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03887_ _03910_ _03892_ _03856_ _03912_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_86_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09794_ _01762_ _04732_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ _03858_ _03188_ _03828_ _03702_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_73_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05957_ _00940_ stack\[7\]\[4\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10278__A2 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ _03208_ _03805_ _03801_ net144 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05888_ stack\[12\]\[6\] stack\[13\]\[6\] _01412_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__B2 mem.mem_dff.code_mem\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ _02867_ _02916_ _02912_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07558_ _02867_ _02862_ _02858_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06509_ mem.mem_dff.code_mem\[0\]\[2\] _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07489_ _02412_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ _01887_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output193_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_158_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10949__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09159_ _04124_ _04166_ _04164_ stack\[1\]\[2\] _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05209__A2 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10202__A2 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11121_ _00713_ clknet_leaf_178_clock stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06009__I1 stack\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11052_ _00644_ clknet_leaf_25_clock delay_cycles\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08520__I _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10003_ _04691_ _04647_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09108__B1 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07382__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__A3 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08331__B2 mem.mem_dff.code_mem\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10905_ _00497_ clknet_leaf_181_clock stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05812__C _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _00428_ clknet_leaf_189_clock stack\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05240__S1 _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10767_ _00359_ clknet_leaf_31_clock net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09831__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08634__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10698_ _00290_ clknet_leaf_62_clock mem.mem_dff.data_mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08398__A1 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08398__B2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06215__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11104__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10181__B _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09898__A1 _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06860_ _02288_ _02319_ _02069_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_67_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05811_ _01274_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06791_ _02263_ _02260_ _02265_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05384__A1 _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ _03656_ _03676_ _03687_ stack\[29\]\[4\] _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05742_ _01285_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _03628_ _03199_ _01637_ _03630_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_05673_ net133 _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ _02751_ _02746_ _02753_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08392_ net120 _02101_ _03578_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ mem.mem_dff.code_mem\[22\]\[0\] _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09822__A1 _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08625__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05439__A2 stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ _02643_ _02635_ _02646_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _04038_ _04063_ _04064_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06225_ _01723_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08389__A1 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08389__B2 _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06156_ _01689_ _01693_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10196__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07061__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06087_ _01624_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09915_ _04819_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09889__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09889__B2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09846_ _01960_ _04759_ _04772_ _03569_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A1 _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ single_step _04262_ _04474_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06989_ _02358_ _02418_ _02408_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06795__I mem.mem_dff.code_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _03844_ _03829_ _03840_ stack\[8\]\[5\] _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_84_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10621__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output206_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ _03656_ _03778_ _03792_ stack\[4\]\[4\] _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A1 _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05517__I3 stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06875__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10110__I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10621_ _00213_ clknet_leaf_105_clock mem.mem_dff.code_mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10771__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08616__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10552_ _00144_ clknet_leaf_79_clock mem.mem_dff.code_mem\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08515__I _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10483_ _00075_ clknet_leaf_56_clock mem.mem_dff.code_mem\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06035__I _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09041__A2 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07575__B _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11104_ _00696_ clknet_leaf_34_clock net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11035_ _00627_ clknet_leaf_22_clock cycles_per_ms\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09081__I _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06315__B1 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10819_ _00411_ clknet_leaf_170_clock stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09804__A1 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08425__I _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ _01405_ _01552_ _01553_ _01416_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xoutput204 net204 rambus_wb_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput215 net239 rambus_wb_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09032__A2 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput226 net226 rambus_wb_rst_o vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08240__B1 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08791__A1 stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ _02998_ _03171_ _03177_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ _04339_ _04473_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06912_ _02314_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07892_ _03124_ _03116_ _03128_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_106_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ cycles_per_ms\[3\] _04586_ _04590_ cycles_per_ms\[2\] _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06843_ _02294_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06829__B _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09562_ cycles_per_ms\[16\] _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06774_ _02128_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08513_ _03191_ _03674_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_05725_ _01264_ stack\[6\]\[2\] _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10794__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09493_ _01286_ _04449_ _04459_ _04337_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input104_I rambus_wb_dat_i[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _03282_ _03244_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05656_ _01199_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08375_ _03561_ _03562_ _03563_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05587_ _01133_ stack\[3\]\[7\] _01105_ stack\[2\]\[7\] _01134_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07326_ _02631_ _02679_ _02686_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07282__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A2 _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _02630_ _02622_ _02633_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06208_ _01181_ _01734_ _01738_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _02489_ _02576_ _02572_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09023__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07034__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06139_ _01137_ _01671_ _01681_ _01648_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08782__B2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output156_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_1_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09829_ _01727_ _04758_ _04760_ _04761_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10341__A1 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07414__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08837__A2 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ _00196_ clknet_leaf_93_clock mem.mem_dff.code_mem\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09262__A2 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10517__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__A1 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _00127_ clknet_leaf_114_clock mem.mem_dff.code_mem\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06076__A2 _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05823__A2 _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10466_ _00058_ clknet_leaf_85_clock mem.mem_dff.code_mem\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09014__A2 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07025__A1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08368__A4 _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ net148 _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10667__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07576__A2 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__A3 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05587__A1 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05587__B2 stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08525__A1 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11018_ _00610_ clknet_leaf_17_clock cycles_per_ms\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08525__B2 stack\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10332__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07324__I mem.mem_dff.code_mem\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08828__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05510_ _00922_ _01059_ _00920_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06490_ net187 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05441_ _00986_ _00987_ _00991_ _00879_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08160_ _02070_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05372_ _00923_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09253__A2 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07111_ _02515_ _02516_ _02518_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07264__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ mem.io_data_out\[7\] _03243_ _03271_ _03287_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_32_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ mem.mem_dff.code_mem\[13\]\[7\] _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__A2 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08764__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08764__B2 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ _03868_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ mem.mem_dff.data_mem\[6\]\[6\] _03163_ _03160_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09714__I _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07875_ mem.mem_dff.data_mem\[4\]\[4\] _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06826_ _02286_ _02293_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09614_ delay_cycles\[4\] _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07234__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09545_ cycles_per_ms\[21\] _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06757_ _02194_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05750__A1 _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__A2 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05708_ _01244_ _01249_ _01251_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09476_ _04442_ _04444_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06688_ _02182_ _02175_ _02184_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08427_ net113 _03603_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05639_ _01182_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05502__A1 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05353__I1 stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08358_ mem.mem_dff.code_mem\[25\]\[7\] _03340_ _03341_ mem.mem_dff.code_mem\[27\]\[7\]
+ _03546_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09244__A2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _02670_ _02663_ _02673_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ mem.mem_dff.data_mem\[0\]\[4\] _03475_ _03476_ _03480_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_203_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10320_ _03858_ _04209_ _04026_ _03233_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_180_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08204__B1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _05059_ _05072_ _05083_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07409__I mem.mem_dff.code_mem\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__B1 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10182_ net171 _05023_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05959__I3 stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout250 net251 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10314__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_210_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_5_0_clock_I clknet_2_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06297__A2 _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__I2 stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06049__A2 _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10250__B1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08994__A1 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10518_ _00110_ clknet_leaf_112_clock mem.mem_dff.code_mem\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ _00041_ clknet_leaf_68_clock mem.mem_dff.code_mem\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08746__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ _01480_ _01530_ _01533_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08349__I1 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09171__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07660_ _02055_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09710__A3 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06611_ _02121_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07591_ _02892_ _02889_ _02893_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09330_ _01833_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06542_ _02064_ _02052_ _02066_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06893__I _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09474__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09261_ _03908_ _04246_ _04233_ _03733_ _04247_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06473_ mem.mem_dff.cycles\[0\] _01995_ _02006_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05335__I1 _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08212_ mem.mem_dff.code_mem\[1\]\[2\] _03355_ _03405_ mem.mem_dff.code_mem\[16\]\[2\]
+ _03356_ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05496__B1 _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05424_ stack\[31\]\[3\] stack\[28\]\[3\] stack\[29\]\[3\] stack\[30\]\[3\] _00968_
+ _00963_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ _04173_ _04196_ _04198_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10832__CLK clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09226__A2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08143_ mem.mem_dff.code_mem\[9\]\[1\] _02321_ _02876_ mem.mem_dff.code_mem\[28\]\[1\]
+ _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05355_ _00815_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08985__A1 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _03253_ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05286_ _00840_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02358_ _02446_ _02437_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10982__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08737__A1 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06133__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08976_ _04013_ _04027_ _04035_ stack\[0\]\[5\] _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input32_I i_wb_addr[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07927_ _03154_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09162__B2 stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ _03101_ _03018_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09701__A3 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__A2 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06809_ _02160_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07789_ _03041_ _03046_ _03048_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output119_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09528_ delay_cycles\[13\] _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08268__A3 _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07476__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _04423_ _04415_ _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05487__B1 _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05212__I _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08976__B2 stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10303_ stack\[27\]\[2\] _05112_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_12_0_clock_I clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06451__A2 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08728__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10234_ _04205_ _05067_ _05070_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06978__I _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _05017_ _05018_ _05010_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10096_ _04949_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08900__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__B2 stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09303__B _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10855__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _00590_ clknet_leaf_129_clock exec.memory_input\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07602__I _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07467__A1 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_9_0_clock_I clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10223__B1 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08967__B2 stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08433__I _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06442__A2 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07049__I _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08719__A1 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09767__I0 exec.memory_input\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08830_ _03924_ _03925_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09264__I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_191_clock clknet_4_0_0_clock clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _03752_ _03864_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05973_ _01426_ _01515_ _01516_ _01430_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05953__A1 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09144__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07712_ _00764_ _01173_ _01174_ _02987_ _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_6_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08692_ _03692_ _03796_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07643_ _02852_ _02931_ _02923_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07574_ mem.mem_dff.code_mem\[28\]\[1\] _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ mem.io_data_out\[2\] _04274_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07458__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ _02051_ _02052_ _02046_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08655__B1 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _04185_ _04235_ _04232_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_179_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06456_ net152 _01716_ _01830_ stack\[2\]\[7\] _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_210_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06130__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11010__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05407_ _00772_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09175_ _03936_ _04182_ _04184_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06387_ _01893_ _01641_ _01924_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09439__I _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ mem.mem_dff.data_mem\[1\]\[0\] _03016_ _03070_ mem.mem_dff.data_mem\[3\]\[0\]
+ mem.mem_dff.data_mem\[7\]\[0\] _03321_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05338_ _00890_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05316__S0 _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_144_clock clknet_4_5_0_clock clknet_leaf_144_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08057_ mem.io_data_out\[1\] _03244_ _03246_ _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06433__A2 _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05269_ stack\[31\]\[0\] stack\[28\]\[0\] stack\[29\]\[0\] stack\[30\]\[0\] _00822_
+ _00823_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11160__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07008_ _02436_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10728__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09383__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput104 rambus_wb_dat_i[4] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_153_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_159_clock clknet_4_6_0_clock clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06197__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05944__A1 _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _01684_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_154_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10878__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A2 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09902__I _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07697__A1 _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _00513_ clknet_leaf_182_clock stack\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06747__B _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10852_ _00444_ clknet_leaf_173_clock stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__B1 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10783_ _00375_ clknet_leaf_135_clock stack\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06672__A2 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07578__B _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08949__A1 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_79_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07621__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05227__A3 _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06424__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10217_ _05057_ _05055_ _05058_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ net238 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A2 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06501__I _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _04565_ _04996_ _05001_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05935__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05935__B2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10079_ _01700_ _04944_ _04946_ intr\[0\] _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08334__C1 mem.mem_dff.code_mem\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11033__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05988__S _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06310_ _01814_ _01809_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07290_ mem.mem_dff.code_mem\[20\]\[3\] _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_206_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06112__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06241_ _00876_ _01782_ _01735_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_61_clock clknet_4_14_0_clock clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05871__B1 _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06172_ _01638_ _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07612__A1 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_76_clock clknet_4_14_0_clock clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09931_ _04819_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08168__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04468_ _04782_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08707__A4 _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07915__A2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08813_ stack\[6\]\[7\] _03896_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _00757_ _04728_ _04734_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05926__B2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05956_ _01485_ stack\[4\]\[4\] _01467_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08744_ _03634_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08675_ _03800_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05887_ _01426_ _01428_ _01429_ _01430_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07626_ mem.mem_dff.code_mem\[29\]\[6\] _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_14_clock clknet_4_8_0_clock clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07557_ _02522_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08628__B1 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06508_ _02035_ _02029_ _02038_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ mem.mem_dff.code_mem\[26\]\[0\] _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06103__A1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29_clock clknet_4_11_0_clock clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09227_ _04175_ _04217_ _04224_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06439_ _01167_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07851__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08073__I _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09158_ _03712_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output186_I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_80_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10550__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08109_ mem.mem_dff.code_mem\[11\]\[0\] _03299_ _03300_ mem.mem_dff.code_mem\[26\]\[0\]
+ _03304_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07603__A1 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09089_ _01792_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08800__B1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ _00712_ clknet_leaf_178_clock stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _00643_ clknet_leaf_25_clock delay_cycles\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10002_ _03627_ _04878_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06321__I _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05917__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09108__A1 _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09108__B2 stack\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07861__B _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _00496_ clknet_leaf_180_clock stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06342__A1 exec.memory_input\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10835_ _00427_ clknet_leaf_189_clock stack\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08095__A1 mem.mem_dff.code_mem\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10766_ _00358_ clknet_leaf_36_clock net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10697_ _00289_ clknet_leaf_62_clock mem.mem_dff.data_mem\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09898__A2 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _00926_ _01352_ _01353_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06790_ _02264_ _02261_ _02252_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06581__A1 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05741_ _00786_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10423__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08460_ _03629_ _03194_ _03195_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08158__I _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05672_ net134 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07411_ _02752_ _02747_ _02743_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _03575_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07997__I _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07342_ _02696_ _02689_ _02698_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08086__A1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09822__A2 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10573__CLK clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07273_ _02644_ _02636_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_102_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09012_ _04040_ _04044_ _04057_ stack\[25\]\[6\] _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ net9 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06155_ _00699_ _01694_ _01697_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_219_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06850__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10196__A2 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__I single_step vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08621__I _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06086_ _01629_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09338__A1 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09914_ _04807_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06141__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08010__A1 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11079__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _04577_ _04757_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07681__B _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _04721_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06572__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06988_ mem.mem_dff.code_mem\[12\]\[2\] _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09452__I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ _03227_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05939_ stack\[18\]\[4\] stack\[19\]\[4\] stack\[16\]\[4\] stack\[17\]\[4\] _00856_
+ _00793_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09510__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08658_ _03782_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A2 _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ _02852_ _02905_ _02898_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ _01990_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10620_ _00212_ clknet_leaf_105_clock mem.mem_dff.code_mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07700__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10551_ _00143_ clknet_leaf_79_clock mem.mem_dff.code_mem\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10482_ _00074_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06316__I _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05220__I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11103_ _00695_ clknet_leaf_34_clock net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11034_ _00626_ clknet_leaf_33_clock cycles_per_ms\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10446__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08304__A2 _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__A1 _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10596__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06935__B _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08068__A1 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08706__I _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _00410_ clknet_leaf_168_clock stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10749_ _00341_ clknet_leaf_38_clock mem.io_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput205 net205 rambus_wb_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput216 net216 rambus_wb_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput227 net227 rambus_wb_sel_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_182_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08791__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ mem.mem_dff.data_mem\[7\]\[3\] _03172_ _03176_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06911_ mem.mem_dff.code_mem\[10\]\[3\] _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07891_ _03125_ _03117_ _03127_ _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09630_ delay_cycles\[2\] _04589_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08543__A2 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06842_ _02294_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06554__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06773_ mem.mem_dff.code_mem\[6\]\[7\] _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09561_ _04509_ _04493_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10939__CLK clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10211__I _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05724_ _01264_ stack\[4\]\[2\] _01267_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08512_ _03638_ _01703_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09492_ _04439_ _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08443_ _02064_ _03609_ _03615_ _03612_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05655_ _01190_ _01192_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08374_ mem.mem_dff.data_mem\[2\]\[7\] _03327_ _03329_ mem.mem_dff.data_mem\[6\]\[7\]
+ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05586_ _01051_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ _02671_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__A1 _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ _02631_ _02623_ _02632_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06207_ _01732_ _01749_ _01181_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07187_ mem.mem_dff.code_mem\[17\]\[5\] _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09023__A3 _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I i_wb_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06138_ _01255_ _01671_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__A1 mem.mem_dff.code_mem\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06069_ _00805_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10469__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06793__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05840__I0 stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output149_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09731__A1 _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ _04336_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _04711_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_185_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__B2 mem.mem_dff.code_mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09910__I _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05215__I _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10603_ _00195_ clknet_leaf_93_clock mem.mem_dff.code_mem\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09798__A1 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10534_ _00126_ clknet_leaf_113_clock mem.mem_dff.code_mem\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ _00057_ clknet_leaf_70_clock mem.mem_dff.code_mem\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09357__I _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07025__A2 _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _05169_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05587__A2 stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__I0 stack\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _00609_ clknet_leaf_41_clock net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07605__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__A2 _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05440_ _00889_ _00989_ _00990_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08436__I _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__B1 _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07340__I _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05371_ _00883_ _00832_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_202_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07110_ _02485_ _02517_ _02513_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10399__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08090_ net119 _03272_ _03286_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07041_ _02461_ _02456_ _02462_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07496__B _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10611__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08171__I _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A2 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09961__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07567__A3 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10206__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _04047_ _04049_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05822__I0 stack\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07943_ _03005_ _03162_ _03165_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__A1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08516__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07874_ _03111_ _03103_ _03114_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07515__I mem.mem_dff.code_mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09613_ _04556_ _04490_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06825_ _02292_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09544_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11117__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06756_ mem.mem_dff.code_mem\[6\]\[3\] _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05750__A2 _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10087__A1 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05707_ _01193_ _01250_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06687_ _02150_ _02176_ _02183_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09475_ _01767_ _01725_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_24_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05889__I0 stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ _02031_ _03602_ _03604_ _03605_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__B1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05638_ _01181_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05353__I2 stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08357_ _03545_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05569_ _01028_ _01117_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09244__A3 _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07308_ _02644_ _02664_ _02672_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ _03477_ _03478_ _03479_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ _02133_ _02618_ _02586_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_153_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10250_ _04222_ _05074_ _05082_ stack\[14\]\[3\] _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_191_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09952__A1 delay_cycles\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__B2 _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _05029_ _05030_ _05022_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout240 net241 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_219_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout251 net252 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06518__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10314__A2 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07191__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_opt_3_0_clock clknet_4_7_0_clock clknet_opt_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08691__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07160__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05895__I3 stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10634__CLK clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08443__A1 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_149_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10517_ _00109_ clknet_leaf_110_clock mem.mem_dff.code_mem\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10250__B2 stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10448_ _00040_ clknet_leaf_69_clock mem.mem_dff.code_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10002__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10784__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10379_ _04915_ _05174_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__A2 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09710__A4 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06610_ net237 _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07590_ _02835_ _02890_ _02886_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06541_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06472_ mem.mem_dff.cycles\[0\] _01995_ _01996_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09260_ stack\[22\]\[6\] _04238_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08682__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08211_ _02535_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05496__A1 stack\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05423_ _00972_ _00973_ _00974_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09191_ _04124_ _04192_ _04189_ stack\[20\]\[2\] _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05496__B2 stack\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08142_ _03337_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05354_ _00894_ _00905_ _00906_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09631__B1 _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10241__A1 _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _03251_ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08985__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05285_ _00839_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07024_ mem.mem_dff.code_mem\[13\]\[2\] _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08975_ _03959_ _04022_ _04036_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07926_ _02467_ _02989_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input25_I i_wb_addr[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__A1 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06808_ mem.mem_dff.code_mem\[7\]\[6\] _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07788_ _02930_ _03047_ _03039_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06920__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ delay_cycles\[14\] _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_45_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06739_ mem.mem_dff.code_mem\[6\]\[0\] _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10657__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ _02009_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05487__A1 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08409_ net124 _02116_ _03591_ _03592_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__05487__B2 stack\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09389_ _04277_ _04364_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_150_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10232__A1 _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08976__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10302_ _03869_ _05117_ _05119_ _05120_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08728__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _04206_ _05051_ _05062_ stack\[12\]\[7\] _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10164_ _04537_ _05008_ _05013_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _04376_ _04961_ _04944_ _01114_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05714__A2 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__C _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10997_ _00589_ clknet_leaf_12_clock edge_interrupts vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__B _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__A1 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10223__B2 stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05650__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09767__I1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ stack\[11\]\[1\] _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05972_ stack\[24\]\[5\] stack\[25\]\[5\] _01374_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05953__A2 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07711_ _02345_ net186 _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08691_ _03794_ _03808_ _03815_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07642_ mem.mem_dff.code_mem\[30\]\[1\] _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07573_ _02873_ _02878_ _02880_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ _04268_ mem.dff_data_out\[2\] _04294_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06524_ _02028_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08655__A1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09852__B1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10057__A4 _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05469__A1 _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09243_ _04235_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06455_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05406_ _00950_ _00957_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08670__A4 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09174_ _03937_ _04162_ _04178_ stack\[1\]\[7\] _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06386_ stack\[2\]\[5\] _01830_ _01923_ _01714_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10214__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08125_ _03320_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05337_ _00767_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09080__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05469__B _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05316__S1 _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08056_ net113 _03250_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05268_ _00802_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07007_ _02376_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07684__B _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05199_ _00758_ net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07394__A1 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput105 rambus_wb_dat_i[5] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08958_ _01757_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05944__A2 stack\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09135__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output131_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ _03112_ _03134_ _03141_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output229_I net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07146__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ _03827_ _03673_ _03944_ _03945_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10920_ _00512_ clknet_leaf_180_clock stack\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__I mem.mem_dff.code_mem\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _00443_ clknet_leaf_0_clock stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10782_ _00374_ clknet_leaf_135_clock stack\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05223__I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__A1 stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08949__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10216_ _04220_ _05050_ _05048_ stack\[12\]\[2\] _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11196_ net241 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ net162 _04999_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10822__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09126__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10078_ _04922_ _04925_ _04945_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08334__C2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A1 stack\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__CLK clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08098__C1 mem.mem_dff.code_mem\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06112__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _01771_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06171_ _01677_ _01685_ _01692_ _01713_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__B2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__B _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _04829_ _04831_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06899__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04551_ _04769_ _04780_ net46 _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _03908_ _03910_ _03892_ _03733_ _03911_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__B _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09792_ net128 _04730_ _04731_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05926__A2 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05482__S0 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ _03854_ _03850_ _03825_ _03856_ _03857_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05955_ _00940_ stack\[5\]\[4\] _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08674_ stack\[5\]\[0\] _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05886_ _01285_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__I _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07625_ _02918_ _02915_ _02919_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06351__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07556_ mem.mem_dff.code_mem\[27\]\[6\] _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08628__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08628__B2 stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06507_ _02037_ _02032_ _02033_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07300__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07487_ _02809_ _02802_ _02811_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06103__A2 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input92_I rambus_wb_dat_i[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09226_ _04222_ _04215_ _04223_ stack\[21\]\[3\] _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06438_ _01780_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05862__A1 _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05862__B2 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09157_ _04169_ _04171_ _04172_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06369_ _01025_ _01868_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_23_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ _03301_ _03302_ _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08261__C1 mem.mem_dff.code_mem\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ _04066_ _04115_ _04121_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08800__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output179_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08039_ _03242_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10845__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06602__I mem.mem_dff.code_mem\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ _00642_ clknet_leaf_25_clock delay_cycles\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07367__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ wb_write_ack _04354_ _01628_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10371__B1 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05917__A2 _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05218__I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09108__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08529__I _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _00495_ clknet_leaf_147_clock stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06342__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _00426_ clknet_leaf_177_clock stack\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08619__A1 stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__B1 _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10765_ _00357_ clknet_leaf_37_clock net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09292__A1 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_190_clock clknet_4_1_0_clock clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_201_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10696_ _00288_ clknet_leaf_59_clock mem.mem_dff.data_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08252__C1 mem.mem_dff.data_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05605__A1 _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09095__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07608__I mem.mem_dff.code_mem\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__B1 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11179_ net242 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06030__A1 _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11000__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06581__A2 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05384__A3 _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05740_ stack\[8\]\[2\] stack\[9\]\[2\] _00857_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A1 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10114__B1 _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_143_clock clknet_4_5_0_clock clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05671_ _01185_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _02522_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11150__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08390_ _03572_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02644_ _02690_ _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10718__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07499__B _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05798__I _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06097__A1 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_158_clock clknet_4_7_0_clock clknet_leaf_158_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08174__I _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ _02614_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _04015_ _03964_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06223_ _01721_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10868__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06154_ _01660_ _01696_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06085_ _01625_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _04816_ _04818_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _01896_ _04759_ _04771_ _03569_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08010__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ exec.memory_input\[7\] _04353_ _04711_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06987_ _02420_ _02417_ _02421_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08726_ _03791_ _03825_ _03843_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05938_ _01471_ _01481_ _01446_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08849__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A3 _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ _01860_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05869_ stack\[24\]\[6\] stack\[25\]\[6\] _01412_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06324__A2 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07608_ mem.mem_dff.code_mem\[29\]\[1\] _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05532__B1 _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08588_ _03732_ _03704_ _03735_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07539_ _02851_ _02848_ _02853_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09274__A1 _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06088__A1 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _00142_ clknet_leaf_76_clock mem.mem_dff.code_mem\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08084__I _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05501__I _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09209_ _04145_ _04209_ _03777_ _03690_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09026__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10481_ _00073_ clknet_leaf_114_clock mem.mem_dff.code_mem\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11102_ _00694_ clknet_leaf_35_clock net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11023__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _00625_ clknet_leaf_19_clock cycles_per_ms\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06012__A1 _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05446__S0 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_clock clknet_4_14_0_clock clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07760__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08259__I _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08304__A3 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__A2 _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06315__A2 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_clock clknet_4_14_0_clock clknet_leaf_75_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_177_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _00409_ clknet_leaf_162_clock stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10748_ _00340_ clknet_leaf_38_clock mem.io_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05411__I _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10679_ _00271_ clknet_leaf_51_clock mem.mem_dff.data_mem\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput206 net206 rambus_wb_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput217 net236 rambus_wb_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput228 net228 rambus_wb_sel_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A2 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clock clknet_4_8_0_clock clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06910_ _02356_ _02349_ _02359_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07890_ _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10335__B1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06003__A1 _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06003__B2 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06841_ mem.mem_dff.code_mem\[8\]\[4\] _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09740__A2 _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _04495_ _04515_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08169__I _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06772_ _02248_ _02241_ _02249_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08511_ _03187_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05723_ _01266_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09491_ _04388_ _01598_ _04457_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07503__A1 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08442_ net119 _03610_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05654_ _01196_ _01197_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ mem.mem_dff.data_mem\[4\]\[7\] _03323_ _03324_ mem.mem_dff.data_mem\[5\]\[7\]
+ _03325_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09256__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05585_ _01093_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07324_ mem.mem_dff.code_mem\[21\]\[3\] _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10690__CLK clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07022__B _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05321__I _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07255_ _02614_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07957__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06206_ _01202_ _01245_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_178_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07186_ _02574_ _02575_ _02577_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11046__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__B1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _01679_ _01650_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input55_I i_wb_data[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06068_ _01093_ _01080_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08788__B _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05840__I1 stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _04629_ _04759_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06545__A2 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _01644_ _04387_ _04254_ _04686_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_39_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ _03820_ _03823_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output211_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _04648_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _00194_ clknet_leaf_103_clock mem.mem_dff.code_mem\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06327__I _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05231__I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _00125_ clknet_leaf_124_clock mem.mem_dff.code_mem\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06481__A1 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ _00056_ clknet_leaf_85_clock mem.mem_dff.code_mem\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08222__A2 _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10395_ _03224_ _05183_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10413__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A1 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06062__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07981__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05831__I1 stack\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _00608_ clknet_leaf_127_clock net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_211_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09722__A2 _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10563__CLK clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05834__C _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07733__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09306__C _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_145_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09238__A1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05370_ _00921_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11069__CLK clknet_opt_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07040_ _02404_ _02457_ _02453_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08452__I _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08213__A2 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _03918_ _04048_ _04044_ _03866_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ mem.mem_dff.data_mem\[6\]\[5\] _03163_ _03160_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05822__I1 stack\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09283__I _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09174__B1 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09713__A2 _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ _03112_ _03104_ _03113_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09612_ cycles_per_ms\[7\] _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06824_ _02288_ _02291_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09543_ _04497_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06755_ _02234_ _02228_ _02236_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09477__A1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06856__B _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05706_ _01224_ _01208_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09474_ _01724_ net43 _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06686_ _02129_ _02183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08425_ _02009_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05889__I1 stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05637_ _00839_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09229__B2 stack\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05353__I3 stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ mem.mem_dff.code_mem\[10\]\[7\] _03343_ _03344_ mem.mem_dff.code_mem\[24\]\[7\]
+ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05568_ _01036_ stack\[19\]\[6\] _01033_ stack\[18\]\[6\] _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07307_ _02671_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ mem.mem_dff.data_mem\[4\]\[4\] net227 _03329_ mem.mem_dff.data_mem\[6\]\[4\]
+ _03381_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05499_ _00933_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09458__I _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07238_ _00760_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ _02563_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08204__A2 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output161_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10011__A2 _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10180_ _04517_ _05020_ _05025_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09952__A2 _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10586__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout241 net214 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout252 net210 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05226__I _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09921__I _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__A2 _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ _00108_ clknet_leaf_110_clock mem.mem_dff.code_mem\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10250__A2 _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_71_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10447_ _00039_ clknet_leaf_69_clock mem.mem_dff.code_mem\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _05169_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07954__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__B1 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A1 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06540_ _02008_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06471_ _02004_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08682__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10459__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08210_ mem.mem_dff.code_mem\[2\]\[2\] _02098_ _02588_ mem.mem_dff.code_mem\[18\]\[2\]
+ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05496__A2 _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05422_ _00878_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09190_ _04169_ _04196_ _04197_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ mem.dff_data_out\[0\] _03333_ _03336_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05353_ stack\[15\]\[2\] stack\[12\]\[2\] stack\[13\]\[2\] stack\[14\]\[2\] _00843_
+ _00891_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08182__I _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08072_ _03249_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10241__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08985__A3 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05284_ _00838_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07023_ _02448_ _02445_ _02449_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06748__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07945__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ _04011_ _04027_ _04035_ stack\[0\]\[4\] _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07925_ _03151_ _03144_ _03153_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07856_ _03098_ _03099_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06807_ _02276_ _02273_ _02277_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input18_I i_wb_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _03045_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09526_ delay_cycles\[15\] _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06738_ _02220_ _02213_ _02222_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_213_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09457_ _04403_ _04427_ _04364_ _04346_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06669_ _02017_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09870__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _03575_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05487__A2 stack\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ _04364_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08339_ _03525_ _03526_ _03527_ _03528_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_178_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06605__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06987__A2 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10301_ _03752_ _05114_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09916__I _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10232_ _05066_ _05067_ _05069_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10163_ net166 _05011_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _04938_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10601__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10996_ _00588_ clknet_leaf_8_clock intr_enable\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__B1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A1 _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__B2 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10751__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10223__A2 _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11107__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08730__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__B1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06250__I _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05971_ stack\[26\]\[5\] stack\[27\]\[5\] _01360_ _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07710_ _02021_ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _03659_ _03800_ _03813_ stack\[5\]\[5\] _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08378__S _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07641_ _02925_ _02929_ _02932_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07572_ _02818_ _02879_ _02871_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07081__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09311_ _04290_ _04293_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06523_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__A1 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08655__A2 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09852__B2 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06666__A1 _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05469__A2 _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ _04145_ _04209_ _03828_ _01712_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_167_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09510__B _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06454_ _01989_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05405_ _00922_ _00952_ _00956_ _00908_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09173_ _04133_ _04182_ _04183_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06385_ _01922_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ _03098_ _02135_ _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06418__A1 _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10214__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05336_ _00887_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07091__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08055_ net70 _03252_ _03254_ net121 _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05267_ _00821_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ mem.mem_dff.code_mem\[12\]\[7\] _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05198_ _00756_ _00757_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput106 rambus_wb_dat_i[6] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08591__A1 _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _04022_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07908_ _03126_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10624__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08888_ _03969_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09471__I _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07839_ _03071_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output124_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10150__A1 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10850_ _00442_ clknet_leaf_169_clock stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09509_ _02004_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10774__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _00373_ clknet_leaf_135_clock stack\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09843__A1 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A2 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__A2 _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__A2 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _03712_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11195_ net242 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10146_ _05003_ _05004_ _04472_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05396__A1 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10077_ net37 _04917_ _04918_ _04931_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08885__A2 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06896__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05699__A2 _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__C1 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10979_ _00571_ clknet_leaf_44_clock net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09834__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05871__A2 _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06170_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09062__A2 _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08270__B1 _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06120__I0 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09860_ _04468_ _04781_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08022__B1 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10647__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08573__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ stack\[6\]\[6\] _03896_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09791_ _03889_ _04732_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10380__A1 _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ stack\[8\]\[7\] _03833_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05482__S1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05954_ _01490_ _01497_ _01424_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08325__A1 mem.mem_dff.code_mem\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08325__B2 mem.mem_dff.code_mem\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08673_ _03802_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10132__A1 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ stack\[8\]\[6\] stack\[9\]\[6\] _01403_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10132__B2 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_193_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07624_ _02835_ _02916_ _02912_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10230__I _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07025__B _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05324__I _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08089__B1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _02864_ _02861_ _02865_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08628__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06506_ _02036_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07486_ _02755_ _02803_ _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _04212_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06437_ _01967_ _01946_ _01971_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input85_I rambus_wb_dat_i[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ _04122_ _04166_ _04164_ stack\[1\]\[1\] _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06368_ _01528_ _01542_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10199__A1 _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09053__A2 _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ mem.mem_dff.code_mem\[25\]\[0\] _02788_ _02845_ mem.mem_dff.code_mem\[27\]\[0\]
+ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05319_ _00864_ _00866_ _00780_ _00872_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09087_ _04024_ _04117_ _04120_ stack\[24\]\[0\] _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08800__A2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06299_ _01803_ _01806_ _01838_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08038_ _03241_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08013__B1 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10000_ _03009_ _04869_ _04877_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05378__A1 _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09989_ _02041_ _04867_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__A1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10371__B2 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05943__B _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10902_ _00494_ clknet_leaf_148_clock stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05925__I0 stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _00425_ clknet_leaf_154_clock stack\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05550__A1 stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08619__A2 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10764_ _00356_ clknet_leaf_37_clock net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09292__A2 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10695_ _00287_ clknet_leaf_62_clock mem.mem_dff.data_mem\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09044__A2 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09376__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05409__I _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__A1 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__B2 _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11178_ net244 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10362__A1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10129_ _04423_ _04961_ _04986_ _04577_ _04140_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05853__B _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06030__A2 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08858__A2 _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__B1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10114__B2 edge_interrupts vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05670_ _01184_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ _02671_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07271_ _02526_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06097__A2 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09010_ _04061_ _04051_ _04062_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06222_ _01763_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09035__A2 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06153_ _01695_ _01658_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08794__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06084_ _01626_ net16 _01627_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_172_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09912_ delay_cycles\[3\] _04811_ _04808_ _04817_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10225__I _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _04592_ _04762_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06986_ _02389_ _02418_ _02408_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09774_ _04344_ _04712_ _04720_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08725_ _03842_ _03829_ _03840_ stack\[8\]\[4\] _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05937_ _01291_ _01475_ _01479_ _01480_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10105__A1 _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _03789_ _03775_ _03790_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__A4 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05907__I0 stack\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _00809_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_215_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07607_ _02900_ _02904_ _02906_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05532__A1 stack\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ stack\[31\]\[6\] _03727_ _03734_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05799_ stack\[2\]\[0\] stack\[3\]\[0\] stack\[0\]\[0\] stack\[1\]\[0\] _00790_ _00802_
+ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05532__B2 stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07538_ _02852_ _02849_ _02842_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09274__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__I1 _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ mem.mem_dff.code_mem\[25\]\[3\] _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09208_ _03187_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10480_ _00072_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10812__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09026__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07037__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09139_ stack\[18\]\[6\] _04149_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07709__I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A1 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05599__A1 _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _00693_ clknet_leaf_33_clock net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__I _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05229__I _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__A1 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _00624_ clknet_leaf_19_clock cycles_per_ms\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10344__A1 _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05446__S1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_9_clock clknet_4_2_0_clock clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08304__A4 _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10816_ _00408_ clknet_leaf_162_clock stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10747_ _00339_ clknet_leaf_38_clock mem.io_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__CLK clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10678_ _00270_ clknet_4_9_0_clock mem.mem_dff.data_mem\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09017__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_141_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07619__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07579__A2 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 net207 rambus_wb_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08776__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06523__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__B1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput218 net234 rambus_wb_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput229 net229 rambus_wb_sel_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A1 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10335__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06840_ _02302_ _02295_ _02304_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09740__A3 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07751__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06771_ _02161_ _02243_ _02238_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08510_ _01675_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05722_ _01265_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09490_ _04442_ _01595_ _04456_ _04387_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_66_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _02060_ _03609_ _03614_ _03612_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05653_ net158 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ mem.mem_dff.data_mem\[1\]\[7\] _03377_ _03378_ mem.mem_dff.data_mem\[3\]\[7\]
+ mem.mem_dff.data_mem\[7\]\[7\] _03321_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10835__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05584_ _01130_ stack\[0\]\[7\] stack\[1\]\[7\] _01131_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09256__A2 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05602__I _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07323_ _02683_ _02678_ _02684_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07254_ _02511_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07019__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06205_ _01635_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07185_ _02485_ _02576_ _02572_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__B2 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06136_ _01652_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_219_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06242__A2 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06067_ _01582_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08519__A1 _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05450__B1 stack\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input48_I i_wb_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09192__A1 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09826_ _04757_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ _04312_ _04475_ _04710_ _04708_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__05753__A1 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06969_ mem.mem_dff.code_mem\[11\]\[7\] _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ _03829_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _04647_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09495__A2 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output204_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _01929_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07213__B _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09247__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10601_ _00193_ clknet_leaf_100_clock mem.mem_dff.code_mem\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09919__I _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10532_ _00124_ clknet_leaf_124_clock mem.mem_dff.code_mem\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _00055_ clknet_leaf_85_clock mem.mem_dff.code_mem\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08758__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ stack\[15\]\[4\] _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08222__A3 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_142_clock clknet_4_5_0_clock clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11140__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10317__A1 _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10708__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _00607_ clknet_leaf_127_clock net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_157_clock clknet_4_7_0_clock clknet_leaf_157_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07733__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06011__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09486__A2 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_202_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05275__A3 _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07349__I _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07421__A1 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04043_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07941_ _03001_ _03162_ _03164_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05983__A1 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09174__B2 stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07872_ _03065_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08921__A1 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _04539_ _04549_ _04553_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06823_ net254 _02290_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06754_ _02235_ _02230_ _02221_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09542_ delay_cycles\[20\] _04496_ delay_cycles\[21\] _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07812__I _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _01246_ _01247_ _01248_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06685_ mem.mem_dff.code_mem\[4\]\[3\] _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08685__B1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _01667_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input102_I rambus_wb_dat_i[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08424_ net112 _03603_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05636_ _01180_ net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09229__A2 _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11013__CLK clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ mem.mem_dff.code_mem\[8\]\[7\] _03292_ _03293_ mem.mem_dff.code_mem\[22\]\[7\]
+ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07968__B _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05567_ _01094_ _01115_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07306_ _02613_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ mem.mem_dff.data_mem\[1\]\[4\] _03016_ _03070_ mem.mem_dff.data_mem\[3\]\[4\]
+ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08643__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05498_ _01042_ stack\[28\]\[5\] stack\[29\]\[5\] _01043_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07237_ mem.mem_dff.code_mem\[19\]\[0\] _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11163__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07168_ _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06119_ net36 net5 _01625_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07099_ _02478_ _02502_ _02495_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_74_clock clknet_4_14_0_clock clknet_leaf_74_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output154_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09407__C _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout242 net243 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout253 net232 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09809_ _02760_ _04744_ _04746_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05726__A1 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_89_clock clknet_4_15_0_clock clknet_leaf_89_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07722__I _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__B1 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_12_clock clknet_4_2_0_clock clknet_leaf_12_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05242__I _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07878__B _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08979__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08553__I _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07651__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _00107_ clknet_leaf_110_clock mem.mem_dff.code_mem\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10446_ _00038_ clknet_leaf_68_clock mem.mem_dff.code_mem\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10530__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06206__A2 _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _03633_ _05172_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08221__C _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__B2 stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10680__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05417__I _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__A2 _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _02003_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05421_ stack\[27\]\[3\] stack\[24\]\[3\] stack\[25\]\[3\] stack\[26\]\[3\] _00968_
+ _00963_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07788__B _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05740__I1 stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08140_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10226__B1 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05352_ _00826_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08463__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__A2 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08071_ _03245_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05283_ _00781_ _00818_ _00837_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08985__A4 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07022_ _02389_ _02446_ _02437_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09395__A1 _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__A2 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06711__I _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _04029_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07924_ _03125_ _03145_ _03152_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05327__I _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07855_ _02289_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05708__A1 _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06806_ _02246_ _02274_ _02270_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07786_ _03045_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ delay_cycles\[18\] _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06737_ _02165_ _02214_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06668_ mem.mem_dff.code_mem\[4\]\[0\] _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _04371_ _04425_ _04426_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08407_ _03572_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05619_ _01126_ _01149_ _01166_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07881__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06599_ _02065_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09387_ _04363_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ mem.mem_dff.code_mem\[17\]\[6\] _03358_ _02620_ mem.mem_dff.code_mem\[19\]\[6\]
+ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08306__C _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ mem.mem_dff.code_mem\[11\]\[4\] _02383_ _02815_ mem.mem_dff.code_mem\[26\]\[4\]
+ _03460_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ stack\[27\]\[1\] _05118_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_188_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09386__A1 _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _05068_ _05051_ _05062_ stack\[12\]\[6\] _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_195_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06621__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _05015_ _05016_ _05010_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10093_ single_step _04941_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05237__I _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__B1 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08361__A2 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08649__B1 _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10995_ _00587_ clknet_leaf_7_clock intr_enable\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09310__A1 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09310__B2 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06124__A1 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__A2 _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10208__B1 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08283__I _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07624__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A1 _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _00021_ clknet_leaf_61_clock mem.mem_dff.code_mem\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05938__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__B2 stack\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05970_ _01462_ _01482_ _01498_ _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09144__A4 _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07640_ _02930_ _02931_ _02923_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10426__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07571_ _02877_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06522_ net241 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09310_ net87 _04291_ _04292_ net79 _04270_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_146_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__A2 _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10576__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09241_ _04233_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06453_ _01983_ _01985_ _01988_ _01649_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05404_ _00894_ _00905_ _00955_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09172_ _04135_ _04162_ _04178_ stack\[1\]\[6\] _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09065__B1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06384_ _01921_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09604__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08123_ _02988_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05335_ _00885_ _00886_ _00887_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10228__I _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__B1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08054_ _02005_ _03257_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05266_ _00820_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _02433_ _02428_ _02434_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05197_ mem.addr\[0\] _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07537__I _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07918__A2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput107 rambus_wb_dat_i[7] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08591__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04021_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input30_I i_wb_addr[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09752__I _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07907_ mem.mem_dff.data_mem\[5\]\[3\] _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08887_ _01640_ _03824_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07838_ _02050_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07272__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07769_ _02943_ _03032_ _03028_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output117_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10919__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ exec.out_of_order_exec _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06106__A1 _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10780_ _00372_ clknet_leaf_10_clock intr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ _01624_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09420__C _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07606__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10138__I _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_197_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__I _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10214_ _05053_ _05055_ _05056_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11194_ net246 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10145_ _04559_ _04996_ _05001_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10449__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10076_ _04943_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06345__A1 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07182__I mem.mem_dff.code_mem\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10599__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08098__A1 mem.mem_dff.code_mem\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__B1 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09295__C2 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10978_ _00570_ clknet_leaf_43_clock net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05430__I _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08270__A1 mem.mem_dff.code_mem\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08741__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08270__B2 mem.mem_dff.code_mem\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06120__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08022__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08022__B2 stack\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _03909_ _03796_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08573__A2 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _04729_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05387__A2 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10380__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _03855_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05953_ _01342_ _01493_ _01496_ _01422_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05884_ stack\[10\]\[6\] stack\[11\]\[6\] _01427_ _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08672_ _03781_ _03800_ _03801_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10132__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ mem.mem_dff.code_mem\[29\]\[5\] _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05934__I1 stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A1 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08089__B2 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ _02835_ _02862_ _02858_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ net248 _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07485_ _02783_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ _01856_ _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06436_ _01967_ _01946_ _01971_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_167_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09589__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ _04170_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06367_ _01900_ _01903_ _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__A2 _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08106_ mem.mem_dff.code_mem\[10\]\[0\] _02346_ _02761_ mem.mem_dff.code_mem\[24\]\[0\]
+ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05318_ _00798_ _00867_ _00871_ _00816_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_175_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I rambus_wb_dat_i[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08651__I _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08261__B2 mem.mem_dff.code_mem\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09086_ _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06298_ _01728_ _01804_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08037_ _00763_ _01177_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05249_ stack\[7\]\[0\] stack\[4\]\[0\] stack\[5\]\[0\] stack\[6\]\[0\] _00801_ _00803_
+ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_150_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__A1 _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__B2 stack\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05378__A2 _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _02994_ _04869_ _04871_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08939_ _04008_ _04001_ _04009_ stack\[13\]\[3\] _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__A2 _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _00493_ clknet_leaf_147_clock stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05925__I1 stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10832_ _00424_ clknet_leaf_153_clock stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10891__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09816__A2 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05550__A2 _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10763_ _00355_ clknet_leaf_37_clock net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09029__B1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _00286_ clknet_4_14_0_clock mem.mem_dff.data_mem\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05250__I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__B _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09044__A3 _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__B2 mem.mem_dff.data_mem\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06081__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09201__B1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06015__B1 _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06566__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ net247 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10362__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ net181 _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__C _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10059_ _04921_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06318__B2 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06030__B _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__B1 _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ mem.mem_dff.code_mem\[19\]\[7\] _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__I _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06221_ _01762_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10614__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06152_ _01657_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_62_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10050__A1 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06083_ net42 net67 _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08794__A2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07087__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09911_ _04586_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10764__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09743__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09842_ _04325_ _04767_ _04770_ _02010_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06557__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09773_ exec.memory_input\[6\] _04712_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ mem.mem_dff.code_mem\[12\]\[1\] _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08724_ _03223_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05936_ _01274_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_4_14_0_clock clknet_3_7_0_clock clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A3 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08655_ _03654_ _03779_ _03783_ stack\[4\]\[3\] _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05867_ stack\[26\]\[6\] stack\[27\]\[6\] _01410_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06875__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05907__I1 stack\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07606_ _02818_ _02905_ _02898_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _03733_ _03717_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05532__A2 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05798_ _01290_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07809__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ _02505_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ _02796_ _02791_ _02797_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__A1 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__B2 stack\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09207_ _03989_ _04087_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_155_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06419_ _01947_ _01954_ _01955_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07399_ _02742_ _02734_ _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__I _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09138_ _03909_ _03662_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output184_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ _03879_ _04095_ _04105_ _04106_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11100_ _00692_ clknet_leaf_35_clock net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__A2 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11031_ _00623_ clknet_4_8_0_clock cycles_per_ms\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05954__B _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06548__A1 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07725__I _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10151__I _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05245__I _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06020__I0 stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08556__I stack\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10815_ _00407_ clknet_leaf_159_clock stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10100__B _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10637__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10746_ _00338_ clknet_leaf_3_clock stack\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10280__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10677_ _00269_ clknet_leaf_49_clock mem.mem_dff.data_mem\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_199_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09387__I _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08291__I _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10787__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net208 rambus_wb_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08776__A2 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput219 net219 rambus_wb_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_141_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09725__A1 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08528__A2 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10335__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__A4 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06770_ mem.mem_dff.code_mem\[6\]\[6\] _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09850__I _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10099__A1 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05721_ _00774_ _00766_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08440_ net118 _03610_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08466__I _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05652_ net258 _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07370__I _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08371_ mem.mem_dff.code_mem\[0\]\[7\] _03451_ _03550_ _03559_ _03473_ _03560_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05583_ _01084_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _02597_ _02679_ _02672_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ mem.mem_dff.code_mem\[19\]\[3\] _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06204_ exec.memory_input\[0\] _01744_ _01746_ _00877_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07184_ _02563_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07019__A2 _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09964__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01598_ _01621_ _01615_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__I _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06066_ _01255_ _01583_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05450__A1 _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__A2 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05450__B2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07545__I _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ _04757_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09192__A2 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09756_ edge_interrupts _04474_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06968_ _02403_ _02398_ _02405_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06950__A1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05753__A2 _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08707_ _03827_ _03673_ _03828_ _03192_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__11092__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05919_ _00880_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ net143 _04641_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06002__I0 stack\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _01757_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ _03715_ _03706_ _03719_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10600_ _00192_ clknet_leaf_100_clock mem.mem_dff.code_mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08455__A1 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10531_ _00123_ clknet_leaf_124_clock mem.mem_dff.code_mem\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08207__A1 _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10462_ _00054_ clknet_leaf_71_clock mem.mem_dff.code_mem\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08758__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10393_ _05182_ _05171_ _05184_ _05185_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09935__I _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11014_ _00606_ clknet_leaf_127_clock net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_10_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08143__B1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09891__B1 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10253__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08997__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ _00321_ clknet_leaf_64_clock mem.mem_dff.data_mem\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06534__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A1 _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A2 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__I0 stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07421__A2 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07940_ mem.mem_dff.data_mem\[6\]\[4\] _03163_ _03160_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07365__I _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09174__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ _02044_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07185__A1 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10005__B _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09610_ _04554_ _04558_ _04562_ _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_214_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06822_ net255 _02289_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08921__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10802__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ delay_cycles\[22\] _04497_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05291__S0 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06753_ _02108_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05704_ _01194_ _01201_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09472_ _01667_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06684_ _02180_ _02175_ _02181_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08685__A1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08685__B2 stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ _03601_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05635_ wb_write_ack wb_read_ack _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _03540_ _03541_ _03542_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08437__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09634__B1 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05566_ _01113_ stack\[16\]\[6\] stack\[17\]\[6\] _01114_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ mem.mem_dff.code_mem\[20\]\[7\] _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10244__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ mem.mem_dff.data_mem\[2\]\[4\] _03043_ _03130_ mem.mem_dff.data_mem\[5\]\[4\]
+ mem.mem_dff.data_mem\[7\]\[4\] _03321_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05497_ _01041_ _01044_ _01046_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_clock clknet_4_2_0_clock clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07236_ _02612_ _02603_ _02616_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _02532_ _02562_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input60_I i_wb_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06118_ _01659_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07098_ mem.mem_dff.code_mem\[15\]\[2\] _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05274__I1 stack\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05423__A1 _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06049_ _01087_ _01252_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout243 net213 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout254 net186 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07176__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09808_ _04406_ _04740_ _04741_ _04745_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10482__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05726__A2 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09739_ _04587_ _04603_ _04600_ _04629_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA_clkbuf_leaf_184_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06619__I _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08676__A1 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__B2 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05523__I _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10235__A1 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08979__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10514_ _00106_ clknet_leaf_115_clock mem.mem_dff.code_mem\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06354__I _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05662__A1 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10445_ _00037_ clknet_leaf_68_clock mem.mem_dff.code_mem\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09665__I cycles_per_ms\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _05168_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05414__A1 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06303__B _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10825__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09156__A2 _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07167__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08903__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07913__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__CLK clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09333__C _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06529__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05433__I _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05420_ _00799_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08419__A1 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08744__I _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05351_ _00903_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08070_ _03263_ _03270_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05282_ _00831_ _00836_ _00781_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07021_ mem.mem_dff.code_mem\[13\]\[1\] _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05405__A1 _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08972_ _03957_ _04023_ _04034_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07095__I _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05956__A2 stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ _03126_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ _02020_ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08919__I _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05708__A2 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06805_ mem.mem_dff.code_mem\[7\]\[5\] _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08370__A3 _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07785_ _03044_ _03018_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__B1 _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _04483_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06736_ _02194_ _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07044__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06439__I _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_141_clock clknet_4_7_0_clock clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09455_ _01124_ _04368_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06667_ _02163_ _02154_ _02167_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_197_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06883__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08406_ net124 _03588_ _03589_ _03086_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11130__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05618_ _01126_ _01165_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08654__I _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _04261_ _04362_ _03625_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06598_ mem.mem_dff.code_mem\[2\]\[3\] _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07881__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08337_ mem.mem_dff.code_mem\[1\]\[6\] _03355_ _03405_ mem.mem_dff.code_mem\[16\]\[6\]
+ _03356_ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05549_ _01009_ _01096_ _01097_ _00938_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_156_clock clknet_4_6_0_clock clknet_leaf_156_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08268_ _03457_ _03458_ _03459_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07219_ _02589_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ mem.mem_dff.code_mem\[23\]\[2\] _03391_ _03392_ mem.mem_dff.code_mem\[31\]\[2\]
+ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10848__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _01124_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10161_ _04542_ _05008_ _05013_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09138__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10092_ _01211_ _04935_ _04951_ intr_enable\[1\] _04139_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10998__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08897__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__B2 stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08361__A3 _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06349__I _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A1 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _00586_ clknet_leaf_10_clock intr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_109_clock clknet_4_13_0_clock clknet_leaf_109_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09310__A2 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06793__B _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08564__I stack\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10208__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10208__B2 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10428_ _00020_ clknet_leaf_61_clock mem.mem_dff.code_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06812__I mem.mem_dff.code_mem\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09377__A2 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _01796_ _05152_ _05160_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09129__A2 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11003__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08739__I _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _02877_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06521_ _02028_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09240_ _04232_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06452_ _01765_ _01986_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_181_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_73_clock clknet_4_14_0_clock clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05403_ stack\[15\]\[3\] stack\[12\]\[3\] stack\[13\]\[3\] stack\[14\]\[3\] _00953_
+ _00954_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09171_ _01932_ _03692_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09065__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06383_ _01821_ _01896_ _01919_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09065__B2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06208__B _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ _02986_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05334_ _00788_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08812__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__B2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08053_ mem.io_data_out\[0\] _03244_ _03246_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_88_clock clknet_4_15_0_clock clknet_leaf_88_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05265_ _00768_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07818__I _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _02404_ _02429_ _02425_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05196_ mem.addr\[1\] _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07379__A1 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05338__I _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06051__A1 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08955_ _01617_ _03201_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput108 rambus_wb_dat_i[8] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07906_ _03138_ _03133_ _03139_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ _03887_ _03965_ _03942_ _03856_ _03968_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I i_wb_addr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07837_ _03071_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_26_clock clknet_4_8_0_clock clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07551__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07768_ _03019_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_57_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _03616_ _04444_ _04259_ _04437_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06719_ _02207_ _02202_ _02208_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10520__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__A1 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07699_ mem.mem_dff.code_mem\[31\]\[6\] _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06106__A2 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08384__I _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09438_ _04260_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_213_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09369_ _01218_ _04315_ _04347_ _04337_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09056__A1 stack\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08803__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05468__I1 stack\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09359__A2 _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06632__I _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11026__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10213_ _04218_ _05050_ _05048_ stack\[12\]\[1\] _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ net247 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05248__I _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06042__A1 _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10144_ net184 _04999_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06042__B2 _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__I _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ _04932_ _04926_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07463__I mem.mem_dff.code_mem\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06079__I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05912__S _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__A1 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10977_ _00569_ clknet_leaf_44_clock net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__B2 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05711__I _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05856__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10329__I _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07638__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06281__A1 _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08558__B1 _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08022__A2 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10365__B1 _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08740_ _03737_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05952_ _01476_ _01494_ _01495_ _01420_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07373__I mem.mem_dff.code_mem\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08671_ _03679_ _03772_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10543__CLK clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05883_ _00880_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07622_ _02914_ _02915_ _02917_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05822__S _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07553_ mem.mem_dff.code_mem\[27\]\[5\] _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08089__A2 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09286__A1 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09286__B2 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06504_ mem.mem_dff.code_mem\[0\]\[1\] _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10693__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ mem.mem_dff.code_mem\[25\]\[7\] _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05621__I _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09223_ _04173_ _04217_ _04221_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__I _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06435_ _01167_ _01968_ _01970_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_195_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09038__A1 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09154_ _01618_ _03989_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06366_ _01528_ _01542_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_10_0_clock clknet_3_5_0_clock clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08105_ mem.mem_dff.code_mem\[12\]\[0\] _02413_ _02441_ mem.mem_dff.code_mem\[13\]\[0\]
+ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08797__B1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05317_ _00825_ _00797_ _00870_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_163_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09085_ _04071_ _04116_ _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06297_ _01357_ _01320_ _01836_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06272__A1 _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ _01991_ _03236_ _03240_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput90 rambus_wb_dat_i[20] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05248_ _00802_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06272__B2 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__A1 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08013__A2 _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10356__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09987_ _04870_ _01782_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__A1 _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08938_ _03998_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06401__B _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output227_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _03954_ _03943_ _03956_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10900_ _00492_ clknet_leaf_186_clock stack\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _00423_ clknet_leaf_157_clock stack\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09277__A1 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10762_ _00354_ clknet_leaf_49_clock mem.dff_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06627__I _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05531__I _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09029__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _00285_ clknet_leaf_54_clock mem.mem_dff.data_mem\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09029__B2 stack\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10416__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09201__A1 _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09201__B2 stack\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06015__A1 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05907__S _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06015__B2 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11176_ net249 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10566__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _04987_ _04988_ _04989_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07193__I mem.mem_dff.code_mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06311__B _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04922_ _04925_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06318__A2 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08712__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09268__A1 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07142__B _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05829__A1 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05829__B2 _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06220_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08752__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06151_ _01666_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10050__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06082_ net68 _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09991__A2 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10909__CLK clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09910_ _04798_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10338__B1 _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05817__S _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ _04593_ _04769_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07754__A1 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _04719_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06984_ _02410_ _02417_ _02419_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _03789_ _03826_ _03841_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05935_ _01476_ _01477_ _01478_ _01420_ _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _01828_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08927__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05866_ _00880_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07605_ _02903_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08585_ _01937_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05797_ stack\[6\]\[0\] stack\[7\]\[0\] _00801_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07536_ mem.mem_dff.code_mem\[27\]\[1\] _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ _02710_ _02792_ _02784_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08482__A2 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input90_I rambus_wb_dat_i[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10439__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04205_ _04203_ _04207_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06418_ _01217_ _01820_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07398_ _02726_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09137_ _04061_ _04143_ _04156_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06349_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07278__I _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__A1 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09068_ _03762_ _04092_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output177_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08019_ _01861_ _03213_ _03226_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11030_ _00622_ clknet_leaf_20_clock cycles_per_ms\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09734__A2 _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06548__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08942__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05526__I _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09498__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05508__B1 _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05359__I0 stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__B _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__I _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06020__I1 stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10814_ _00406_ clknet_leaf_161_clock stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _00337_ clknet_leaf_3_clock stack\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06484__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10280__A2 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10676_ _00268_ clknet_leaf_48_clock mem.mem_dff.data_mem\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput209 net209 rambus_wb_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__A2 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_179_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__I _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09725__A2 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__C _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07736__A1 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11159_ _00751_ clknet_leaf_168_clock stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05720_ _01014_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10099__A2 _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05651_ _01189_ _01194_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03551_ _03552_ _03557_ _03558_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05582_ _01083_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07321_ mem.mem_dff.code_mem\[21\]\[2\] _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09578__I _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07252_ _02628_ _02622_ _02629_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06203_ _01745_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10731__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07183_ _02563_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06227__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06134_ _01676_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06065_ _01279_ _01591_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10881__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05450__A2 stack\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09716__A2 _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__A3 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _04756_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05346__I _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06967_ _02404_ _02399_ _02395_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09755_ _03623_ _04706_ _04709_ _04708_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06886__B _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06950__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05918_ _01454_ _01461_ _01424_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08706_ _01929_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09686_ _04253_ _04480_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08657__I _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06898_ net249 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07561__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06002__I1 stack\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08637_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05849_ stack\[6\]\[7\] stack\[7\]\[7\] _01369_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_4_0_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08568_ _03221_ _03711_ _03718_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07519_ mem.mem_dff.code_mem\[26\]\[6\] _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08499_ _03640_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10530_ _00122_ clknet_leaf_112_clock mem.mem_dff.code_mem\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _00053_ clknet_leaf_72_clock mem.mem_dff.code_mem\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08207__A2 _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06218__A1 _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_180_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _04103_ _05174_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06769__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09707__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07981__A4 _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07718__A1 _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11013_ _00605_ clknet_4_12_0_clock net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05256__I _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09891__A1 _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08694__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09891__B2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09900__B _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05752__I0 stack\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05920__S _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10754__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09398__I _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06457__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10728_ _00320_ clknet_leaf_64_clock mem.mem_dff.data_mem\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10253__A2 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10659_ _00251_ clknet_leaf_78_clock mem.mem_dff.code_mem\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06209__A1 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__A2 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07957__A1 mem.mem_dff.data_mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05807__I1 stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07646__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09159__B1 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06550__I _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__B1 _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05983__A3 _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ mem.mem_dff.data_mem\[4\]\[3\] _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A1 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__C _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06821_ _00758_ _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08921__A3 _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09540_ cycles_per_ms\[22\] _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06752_ mem.mem_dff.code_mem\[6\]\[2\] _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05291__S1 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08134__A1 mem.mem_dff.data_mem\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07381__I mem.mem_dff.code_mem\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05991__I0 stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05703_ _01199_ _01201_ _01213_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_184_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _04387_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06683_ _02109_ _02176_ _02166_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08685__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08422_ _03601_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05634_ edge_interrupts prev_level_interrupt _01179_ net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08353_ mem.mem_dff.code_mem\[23\]\[7\] _02730_ _02956_ mem.mem_dff.code_mem\[31\]\[7\]
+ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05565_ _00969_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09634__A1 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09634__B2 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07304_ _02668_ _02663_ _02669_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06448__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10244__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06725__I _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _02988_ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05496_ stack\[26\]\[5\] _01045_ _00960_ stack\[27\]\[5\] _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ _02527_ _02605_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07166_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ net35 net4 _01654_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07097_ _02504_ _02501_ _02507_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input53_I i_wb_data[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05423__A2 _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05274__I2 stack\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _01260_ _01591_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout233 net234 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout244 net245 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10627__CLK clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout255 net185 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09807_ _01859_ _04739_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10180__A1 _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ _03208_ _03209_ _03210_ net144 _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09738_ _04540_ _04537_ _04542_ _04551_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_74_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_127_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10777__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09873__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ cycles_per_ms\[0\] _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08676__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06687__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05740__S _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06635__I mem.mem_dff.code_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _00105_ clknet_leaf_115_clock mem.mem_dff.code_mem\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10157__I _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09946__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10444_ _00036_ clknet_leaf_74_clock mem.mem_dff.code_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08850__I _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05662__A2 _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05695__B _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10375_ _05170_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07466__I mem.mem_dff.code_mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__S _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__B2 mem.mem_dff.code_mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08667__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout240_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10226__A2 _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05350_ stack\[11\]\[2\] stack\[8\]\[2\] stack\[9\]\[2\] stack\[10\]\[2\] _00901_
+ _00902_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10067__I _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05281_ _00819_ _00833_ _00835_ _00807_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07020_ _02439_ _02445_ _02447_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06850__A1 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11082__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07376__I mem.mem_dff.code_mem\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08971_ _04008_ _04028_ _04030_ stack\[0\]\[3\] _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07922_ mem.mem_dff.data_mem\[5\]\[7\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09591__I cycles_per_ms\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08355__B2 mem.mem_dff.code_mem\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07853_ mem.mem_dff.data_mem\[4\]\[0\] _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06804_ _02272_ _02273_ _02275_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08370__A4 _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07784_ _03043_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__A1 mem.mem_dff.code_mem\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06735_ mem.mem_dff.code_mem\[5\]\[7\] _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09523_ cycles_per_ms\[23\] _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09454_ _04423_ _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_213_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06666_ _02165_ _02155_ _02166_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08405_ _03575_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05617_ _01153_ _01157_ _01160_ _01164_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09385_ _04361_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06597_ _02107_ _02100_ _02110_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ mem.mem_dff.code_mem\[2\]\[6\] _02098_ _02588_ mem.mem_dff.code_mem\[18\]\[6\]
+ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10217__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05548_ stack\[6\]\[6\] _01049_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06455__I _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ mem.mem_dff.code_mem\[12\]\[4\] _02413_ _02441_ mem.mem_dff.code_mem\[13\]\[4\]
+ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05479_ _00953_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07218_ mem.mem_dff.code_mem\[18\]\[4\] _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ _02956_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07149_ _02537_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10160_ net165 _05011_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04954_ _04958_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09715__B single_step vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08897__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08361__A4 _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05534__I _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10993_ _00585_ clknet_leaf_13_clock net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09846__A1 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A2 _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08845__I _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10208__A2 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09074__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08282__B1 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06832__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _00019_ clknet_leaf_60_clock mem.mem_dff.code_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _01825_ _05154_ _05157_ stack\[17\]\[2\] _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10392__A1 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10289_ _03186_ _03188_ _03828_ _03702_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08337__B2 mem.mem_dff.code_mem\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10144__A1 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__I _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_clock clknet_4_2_0_clock clknet_leaf_7_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05571__A1 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09837__A1 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06520_ mem.mem_dff.code_mem\[0\]\[4\] _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08755__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06451_ _01765_ net64 _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05402_ _00884_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09170_ _04180_ _04170_ _04181_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06275__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06382_ _01233_ _01737_ _01754_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09065__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08121_ mem.mem_dff.code_mem\[0\]\[0\] _03290_ _03297_ _03315_ _03316_ _03317_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_30_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05333_ stack\[27\]\[2\] stack\[24\]\[2\] stack\[25\]\[2\] stack\[26\]\[2\] _00882_
+ _00884_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_175_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ net112 _03250_ _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06823__A1 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05264_ _00798_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07003_ mem.mem_dff.code_mem\[12\]\[6\] _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09368__A3 _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10383__A1 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06051__A2 _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 rambus_wb_dat_i[9] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_08954_ _04019_ _04017_ _03992_ _03987_ _04020_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_131_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07905_ _03079_ _03134_ _03127_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08885_ stack\[26\]\[7\] _03950_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07836_ mem.mem_dff.data_mem\[3\]\[4\] _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input16_I i_la_wb_disable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ _03019_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05562__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ _01661_ _04259_ _04261_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06718_ _02109_ _02203_ _02195_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07698_ _02975_ _02972_ _02976_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06106__A3 _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06649_ mem.mem_dff.code_mem\[3\]\[4\] _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09437_ _04403_ _04409_ _04399_ _04326_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10815__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__I _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _04264_ _04345_ _04346_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09056__A2 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ mem.mem_dff.data_mem\[0\]\[5\] _03475_ _03476_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09299_ _04268_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08803__A2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05468__I2 stack\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10965__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05529__I _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08567__A1 _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10212_ _05054_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11192_ net251 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10374__A1 _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10143_ _05000_ _05002_ _04472_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10074_ _04258_ _04941_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10126__A1 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09819__A1 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09295__A2 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10976_ _00568_ clknet_leaf_42_clock net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10495__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05856__A2 _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06095__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08558__A1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_140_clock clknet_4_7_0_clock clknet_leaf_140_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10365__A1 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11120__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I i_la_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05951_ stack\[30\]\[4\] stack\[31\]\[4\] _01374_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10117__A1 _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ _03741_ _03637_ _03777_ _03691_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05882_ _01010_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07621_ _02831_ _02916_ _02912_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _02860_ _02861_ _02863_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05902__I _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06503_ _02012_ _02029_ _02034_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07297__A1 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07483_ _02807_ _02802_ _02808_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09222_ _04220_ _04215_ _04213_ stack\[21\]\[2\] _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06434_ _01168_ _01901_ _01867_ _01969_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09038__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ _03868_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10988__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06365_ _01901_ _01902_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07829__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ _02814_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08797__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05316_ stack\[11\]\[1\] stack\[8\]\[1\] stack\[9\]\[1\] stack\[10\]\[1\] _00868_
+ _00869_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_163_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09084_ _03820_ _03940_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06296_ _01357_ _01277_ _01294_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08035_ net152 _03210_ _03225_ stack\[28\]\[7\] _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05247_ _00766_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06272__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput80 rambus_wb_dat_i[11] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput91 rambus_wb_dat_i[21] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08549__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_108_clock clknet_4_13_0_clock clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10356__A1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09986_ _04865_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _01856_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10108__A1 _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05783__A1 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _03837_ _03947_ _03955_ stack\[26\]\[2\] _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07819_ _03070_ _03018_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output122_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08799_ _03895_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10830_ _00422_ clknet_leaf_153_clock stack\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06908__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__A2 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07288__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10761_ _00353_ clknet_leaf_37_clock mem.dff_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10692_ _00284_ clknet_leaf_55_clock mem.mem_dff.data_mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09029__A2 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08788__A1 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09201__A2 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07212__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11175_ clknet_opt_4_1_clock net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_72_clock clknet_4_15_0_clock clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10126_ net180 _04957_ _03183_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10057_ net34 _01655_ _04923_ _04924_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_209_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08712__B2 stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_clock clknet_4_15_0_clock clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_175_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A2 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07279__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10959_ _00551_ clknet_leaf_142_clock stack\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05829__A2 _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_clock clknet_4_3_0_clock clknet_leaf_10_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08228__B1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__A1 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09976__B1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06150_ _00699_ _01668_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06553__I mem.mem_dff.code_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_clock clknet_4_8_0_clock clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_172_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06081_ net17 _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10050__A3 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10338__A1 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10510__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09840_ _04768_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__B _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08951__A1 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ exec.memory_input\[5\] _04333_ _04715_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06983_ _02351_ _02418_ _02408_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _03839_ _03830_ _03840_ stack\[8\]\[3\] _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05934_ stack\[6\]\[3\] stack\[7\]\[3\] _00821_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08703__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05865_ _01010_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08653_ _03787_ _03775_ _03788_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07604_ _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09259__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05796_ stack\[4\]\[0\] stack\[5\]\[0\] _00843_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08584_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11016__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _02844_ _02848_ _02850_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__B1 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07466_ mem.mem_dff.code_mem\[25\]\[2\] _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09205_ _04206_ _04193_ _04200_ stack\[20\]\[7\] _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06417_ _01743_ _01948_ _01953_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _02511_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input83_I rambus_wb_dat_i[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06463__I _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _04131_ _04146_ _04153_ stack\[18\]\[5\] _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06348_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09067_ stack\[23\]\[4\] _04096_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06279_ _01736_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _03224_ _03193_ _03225_ stack\[28\]\[4\] _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09734__A3 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_8_0_clock clknet_3_4_0_clock clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_131_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08942__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08942__B2 stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _04857_ _04858_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09498__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05508__A1 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05359__I1 stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05508__B2 stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _00405_ clknet_leaf_159_clock stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08853__I _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10744_ _00336_ clknet_leaf_170_clock stack\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09670__A2 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07681__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06484__A2 _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10675_ _00267_ clknet_leaf_49_clock mem.mem_dff.data_mem\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06236__A2 _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__B1 _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09725__A3 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10683__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05717__I _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11158_ _00750_ clknet_leaf_133_clock stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10109_ _04968_ _04141_ _04972_ _04974_ _04776_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11089_ _00681_ clknet_leaf_15_clock net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09489__A2 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11039__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05650_ _01191_ _01192_ _01193_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05581_ _01041_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ _02681_ _02678_ _02682_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07251_ _02597_ _02623_ _02615_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ _01247_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ mem.mem_dff.code_mem\[17\]\[4\] _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06283__I _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06133_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06227__A2 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05828__S _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06064_ _01575_ _01232_ _01089_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05986__A1 _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09823_ _01694_ _04362_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_48_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08003__I _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09754_ intr_enable\[1\] _04706_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06966_ _02160_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07842__I mem.mem_dff.data_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ _03634_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05917_ _01408_ _01457_ _01460_ _01422_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09685_ delay_cycles\[23\] _04498_ _04642_ _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__B1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06897_ _02348_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06458__I _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08636_ _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05848_ stack\[4\]\[7\] stack\[5\]\[7\] _01391_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06163__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05910__A1 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _03716_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05779_ stack\[26\]\[0\] stack\[27\]\[0\] _00792_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__B1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _02834_ _02830_ _02836_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _01931_ _03661_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07449_ mem.mem_dff.code_mem\[24\]\[7\] _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _00052_ clknet_leaf_85_clock mem.mem_dff.code_mem\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_123_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09119_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06218__A2 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08612__B1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _03221_ _05183_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09707__A3 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11012_ _00604_ clknet_leaf_127_clock net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05729__A1 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06154__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05272__I _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05901__A1 _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05752__I1 stack\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08583__I _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10727_ _00319_ clknet_leaf_64_clock mem.mem_dff.data_mem\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06457__A2 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10658_ _00250_ clknet_leaf_93_clock mem.mem_dff.code_mem\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _00181_ clknet_leaf_88_clock mem.mem_dff.code_mem\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07927__I _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06831__I mem.mem_dff.code_mem\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__C _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05968__A1 _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__B2 stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__B2 stack\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08382__A2 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06820_ _02287_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10429__CLK clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__A4 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ _02232_ _02228_ _02233_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05702_ _01206_ _01199_ _01201_ _01245_ _01223_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06682_ mem.mem_dff.code_mem\[4\]\[2\] _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09470_ _04438_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06145__A1 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08421_ _02985_ _02256_ _03248_ _03570_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_184_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05633_ intr_enable\[0\] intr\[0\] intr\[1\] intr_enable\[1\] _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08352_ mem.mem_dff.code_mem\[6\]\[7\] _02225_ _02926_ mem.mem_dff.code_mem\[30\]\[7\]
+ _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05564_ _01029_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09634__A2 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07303_ _02641_ _02664_ _02660_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08283_ _02986_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05495_ _00984_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07234_ _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _02069_ _02534_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05259__I0 stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10401__B1 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06116_ _01657_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08070__A1 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07096_ _02506_ _02502_ _02495_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06047_ _01577_ _01322_ _01573_ _01590_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_156_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05274__I3 stack\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I i_wb_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout234 net218 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout245 net246 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout256 net142 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08373__A2 _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _04731_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10180__A2 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _03203_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09737_ cycles_per_ms\[11\] _04565_ _04559_ _04554_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06949_ mem.mem_dff.code_mem\[11\]\[2\] _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ _04597_ _04599_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output202_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08619_ stack\[3\]\[4\] _03760_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09599_ cycles_per_ms\[9\] _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07636__A1 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10512_ _00104_ clknet_leaf_115_clock mem.mem_dff.code_mem\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09389__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10443_ _00035_ clknet_leaf_74_clock mem.mem_dff.code_mem\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06651__I _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10374_ _03261_ _05168_ _05169_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10173__I _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05267__I _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09962__I _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_5_0_clock clknet_2_2_0_clock clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06375__A1 exec.memory_input\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09313__A1 mem.io_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06098__I _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07627__A1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10348__I _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout233_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06047__B _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05280_ _00825_ _00826_ _00834_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06850__A2 _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A1 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08970_ _03954_ _04023_ _04033_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ _03149_ _03144_ _03150_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07852_ _03094_ _03085_ _03096_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07606__B _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06366__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A2 _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06803_ _02242_ _02274_ _02270_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06002__S _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 i_la_addr[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07783_ _02381_ _03042_ _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08107__A2 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09522_ _01171_ _04481_ _04482_ _04467_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06734_ _02218_ _02213_ _02219_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05841__S _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09453_ net155 _04405_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06665_ _02129_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input100_I rambus_wb_dat_i[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08404_ _03572_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05877__B1 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07341__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06736__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05616_ _01162_ _01163_ _01137_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09384_ _01659_ _04360_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06596_ _02109_ _02103_ _02092_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05640__I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08335_ mem.mem_dff.code_mem\[5\]\[6\] _02200_ _02650_ mem.mem_dff.code_mem\[20\]\[6\]
+ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05547_ _01012_ stack\[4\]\[6\] stack\[5\]\[6\] _01043_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08266_ mem.mem_dff.code_mem\[25\]\[4\] _03340_ _03341_ mem.mem_dff.code_mem\[27\]\[4\]
+ _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05478_ _00961_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07217_ _02599_ _02590_ _02601_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08197_ _02730_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06471__I _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ mem.mem_dff.code_mem\[16\]\[4\] _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09791__A1 _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ _02491_ _02484_ _02492_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10090_ net161 _04957_ _04429_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output152_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10744__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06109__A1 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _00584_ clknet_leaf_13_clock net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10894__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06646__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__B1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__B2 _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10426_ _00018_ clknet_leaf_55_clock mem.mem_dff.code_mem\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08034__A1 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09782__A1 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10357_ _03869_ _05152_ _05159_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06596__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10392__A2 _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10288_ _03854_ _05105_ _05108_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07426__B _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06450_ net15 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06556__I mem.mem_dff.code_mem\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05401_ _00926_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06381_ _01729_ _01912_ _01915_ _01918_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_203_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _02015_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10617__CLK clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05332_ stack\[31\]\[2\] stack\[28\]\[2\] stack\[29\]\[2\] stack\[30\]\[2\] _00882_
+ _00884_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08273__A1 mem.mem_dff.code_mem\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ net69 _03252_ _03254_ net120 _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05263_ _00796_ _00808_ _00813_ _00817_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06823__A2 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07002_ _02431_ _02428_ _02432_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06291__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09222__B1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__A2 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__A2 _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ stack\[13\]\[7\] _03999_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07904_ mem.mem_dff.data_mem\[5\]\[2\] _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ _03963_ _03965_ _03966_ _03967_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09107__I _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07835_ _03081_ _03072_ _03083_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08011__I _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ mem.mem_dff.data_mem\[1\]\[4\] _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _04468_ _03570_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06717_ mem.mem_dff.code_mem\[5\]\[2\] _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ _02947_ _02973_ _02969_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07071__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04371_ _04405_ _04407_ _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06648_ _02148_ _02139_ _02152_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _04324_ _01960_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06579_ _02024_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11024__D _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08318_ _03506_ _03507_ _03508_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09298_ net89 _03099_ _04280_ _04281_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _03435_ _03440_ _03441_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05468__I3 stack\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10211_ _05051_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08567__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ net234 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10374__A2 _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _04554_ _04996_ _05001_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput190 net190 rambus_wb_addr_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_95_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10073_ _04933_ _04925_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__A2 _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05545__I _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06750__A1 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11072__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10975_ _00567_ clknet_leaf_45_clock net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_171_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07000__I mem.mem_dff.code_mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09755__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08558__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _00001_ clknet_4_7_0_clock stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06569__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10365__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05950_ stack\[28\]\[4\] stack\[29\]\[4\] _01329_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2_0_clock clknet_0_clock clknet_2_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05881_ _01407_ _01423_ _01424_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _02903_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06741__A1 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05391__S _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07551_ _02831_ _02862_ _02858_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11192__I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_96_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06502_ _02031_ _02032_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05404__B _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07482_ _02752_ _02803_ _02799_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09221_ _01824_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06433_ _01074_ _01122_ _01907_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_50_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09152_ _04165_ _04168_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06364_ _01072_ _01772_ _01899_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_202_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08103_ _02382_ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10053__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09994__A1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05315_ _00784_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08797__A2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _04116_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06295_ _01834_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05855__I0 stack\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08034_ _01964_ _03236_ _03239_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput70 io_in[1] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_135_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05246_ _00800_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput81 rambus_wb_dat_i[12] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput92 rambus_wb_dat_i[22] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_150_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09746__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10356__A2 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _04865_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08936_ _03954_ _04003_ _04007_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10108__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06980__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08867_ _03949_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07818_ _03069_ _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08798_ _03785_ _03901_ _03902_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output115_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07749_ _02014_ _02988_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09277__A3 _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10760_ _00352_ clknet_leaf_48_clock mem.dff_data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08485__A1 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__B2 stack\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05299__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ _04300_ _04384_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_4_0_clock clknet_3_2_0_clock clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_13_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10691_ _00283_ clknet_leaf_59_clock mem.mem_dff.data_mem\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10932__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06924__I _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05968__C _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08788__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_clock clknet_4_2_0_clock clknet_leaf_6_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09737__A1 cycles_per_ms\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05471__A1 _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _01233_ _04969_ _04928_ _01075_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09970__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ net26 net25 net28 net27 _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06023__I0 stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08712__A2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09760__I1 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_118_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08476__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10958_ _00550_ clknet_leaf_141_clock stack\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10283__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10889_ _00481_ clknet_leaf_181_clock stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06834__I mem.mem_dff.code_mem\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05837__I0 stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06080_ net143 _01623_ net141 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10050__A4 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10338__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_217_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08400__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09770_ _04718_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08951__A2 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06982_ _02416_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__CLK clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _03832_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05933_ stack\[4\]\[3\] stack\[5\]\[3\] _01417_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06014__I0 stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08703__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ _03652_ _03779_ _03783_ stack\[4\]\[2\] _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05864_ _01281_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07603_ _02874_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _01962_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10955__CLK clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05795_ _01335_ _01338_ _01321_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06190__A2 _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07534_ _02818_ _02849_ _02842_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10274__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07465_ _02794_ _02791_ _02795_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _01170_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08219__A1 mem.mem_dff.data_mem\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06416_ _01075_ _01780_ _01950_ _01952_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_183_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07396_ mem.mem_dff.code_mem\[23\]\[3\] _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05788__C _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09120__I _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04059_ _04143_ _04155_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06347_ _01821_ _01864_ _01884_ _01885_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_163_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05828__I0 stack\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input76_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09066_ _04102_ _04104_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _01801_ _01807_ _01813_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05453__A1 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09719__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05453__B2 _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08017_ _03204_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05229_ _00775_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08942__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10485__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09968_ delay_cycles\[19\] _04854_ _04852_ _04511_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09790__I _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output232_I net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _03187_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09723__C _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09899_ _04807_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06005__I0 stack\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05508__A2 stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05359__I2 stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _00404_ clknet_leaf_171_clock stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10743_ _00335_ clknet_leaf_167_clock stack\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11110__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06654__I mem.mem_dff.code_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10674_ _00266_ clknet_leaf_59_clock mem.mem_dff.code_mem\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10017__A1 delay_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09958__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10017__B2 _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_154_clock clknet_4_5_0_clock clknet_leaf_154_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10109__C _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08630__A1 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08630__B2 stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_44_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07984__A3 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08090__B _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07485__I _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10828__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_169_clock clknet_4_3_0_clock clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08933__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11157_ _00749_ clknet_leaf_133_clock stack\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05934__S _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10108_ _04100_ _04973_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _00680_ clknet_leaf_128_clock net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10978__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10039_ _04907_ _04908_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05580_ stack\[7\]\[7\] stack\[4\]\[7\] stack\[5\]\[7\] stack\[6\]\[7\] _01113_ _01114_
+ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_107_clock clknet_4_13_0_clock clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10256__A1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ mem.mem_dff.code_mem\[19\]\[2\] _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06564__I _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07672__A2 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06201_ _01246_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07181_ _02571_ _02564_ _02573_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06132_ _01649_ _01651_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05435__A1 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06063_ _01597_ _01606_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07609__B _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05986__A2 _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06005__S _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _04375_ _04440_ _04646_ _04755_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08924__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05294__S0 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09753_ _01727_ _04706_ _04707_ _04708_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06965_ mem.mem_dff.code_mem\[11\]\[6\] _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ _03825_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05916_ _01416_ _01458_ _01459_ _01420_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09684_ _04483_ _04643_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08688__A1 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09885__B1 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ _02286_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__B2 stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08152__A3 _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08635_ _03201_ _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05847_ _00899_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _03699_ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05778_ _01295_ _01320_ _01321_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__A1 _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _02835_ _02832_ _02827_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10247__B2 stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09101__A2 _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03636_ _01925_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07448_ _02780_ _02775_ _02781_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71_clock clknet_4_14_0_clock clknet_leaf_71_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _02644_ _02718_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09118_ _04142_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output182_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08612__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _05168_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08612__B2 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05426__A1 _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_clock clknet_4_15_0_clock clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09049_ stack\[23\]\[0\] _04090_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05977__A2 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11011_ _00603_ clknet_leaf_46_clock net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05729__A2 stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08679__A1 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_clock clknet_4_8_0_clock clknet_leaf_24_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09628__B1 _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05752__I2 stack\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10500__CLK clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10726_ _00318_ clknet_leaf_51_clock mem.mem_dff.data_mem\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_39_clock clknet_4_8_0_clock clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06384__I _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_clock clknet_2_0_0_clock clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_220_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10657_ _00249_ clknet_leaf_95_clock mem.mem_dff.code_mem\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05929__S _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10650__CLK clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ _00180_ clknet_leaf_88_clock mem.mem_dff.code_mem\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07429__B _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05968__A2 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A2 _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08104__I _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08367__B1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__A3 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07590__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06750_ _02144_ _02230_ _02221_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06559__I mem.mem_dff.code_mem\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05463__I _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05701_ _01211_ _01212_ _01235_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09331__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06681_ _02178_ _02175_ _02179_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ _03594_ _03599_ _03600_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05632_ _01178_ net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_184_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_0_0_clock_I clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ mem.mem_dff.code_mem\[15\]\[7\] _02498_ _02901_ mem.mem_dff.code_mem\[29\]\[7\]
+ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05563_ stack\[23\]\[6\] stack\[20\]\[6\] stack\[21\]\[6\] stack\[22\]\[6\] _01030_
+ _01031_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07302_ mem.mem_dff.code_mem\[20\]\[6\] _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08282_ mem.mem_dff.code_mem\[0\]\[4\] _03451_ _03456_ _03472_ _03473_ _03474_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05494_ _01042_ stack\[24\]\[5\] stack\[25\]\[5\] _01043_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08842__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ mem.mem_dff.code_mem\[17\]\[0\] _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05259__I1 stack\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10401__A1 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06115_ net34 net3 net17 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10401__B2 stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07095_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05638__I _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06046_ _01239_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout235 net217 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout246 net212 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I i_wb_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _02813_ _04728_ _04743_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout257 net150 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07997_ _03193_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09736_ _04692_ _04693_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06948_ _02388_ _02385_ _02390_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06469__I _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09667_ _04513_ _04518_ _04523_ _04527_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__10523__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06879_ _02322_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08530__B1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _03745_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09598_ _04555_ _04557_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ _01676_ _03701_ _01691_ _03702_ _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10673__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _00103_ clknet_leaf_115_clock mem.mem_dff.code_mem\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__B _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _00034_ clknet_leaf_68_clock mem.mem_dff.code_mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06932__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11029__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10373_ _03870_ _03991_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09561__A2 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07572__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08116__A3 _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08594__I _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__I mem.mem_dff.code_mem\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10709_ _00301_ clknet_leaf_37_clock mem.mem_dff.data_mem\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08543__B _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07938__I _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06842__I _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09358__C _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ _03122_ _03145_ _03141_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05810__A1 _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08769__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05249__S0 _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _02981_ _03087_ _03095_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10546__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07563__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06802_ _02259_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06289__I _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 i_la_addr[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07782_ _00761_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09521_ _01171_ _04479_ _04481_ _04253_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06733_ _02161_ _02214_ _02210_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06118__A2 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_166_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ net156 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10696__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06664_ _02164_ _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08403_ _03581_ _03586_ _03587_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05877__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05421__S0 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05615_ _01133_ stack\[27\]\[7\] _01140_ stack\[26\]\[7\] _01134_ _01163_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09068__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05877__B2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09383_ _01630_ _03616_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06595_ _02108_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08334_ mem.mem_dff.code_mem\[3\]\[6\] _02137_ _02173_ mem.mem_dff.code_mem\[4\]\[6\]
+ mem.mem_dff.code_mem\[21\]\[6\] _02676_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05546_ _01093_ stack\[3\]\[6\] _01094_ stack\[2\]\[6\] _01051_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ mem.mem_dff.code_mem\[10\]\[4\] _02347_ _02762_ mem.mem_dff.code_mem\[24\]\[4\]
+ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05477_ _01027_ net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07216_ _02512_ _02592_ _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08196_ mem.mem_dff.code_mem\[6\]\[2\] _03388_ _03389_ mem.mem_dff.code_mem\[30\]\[2\]
+ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07147_ _02545_ _02538_ _02547_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__A2 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05368__I _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07078_ _02404_ _02486_ _02481_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05801__A1 _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05801__B2 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06029_ _01359_ _01448_ _01514_ _01572_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_134_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08346__A3 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output145_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07554__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06357__A2 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xspell_260 o_wb_data[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _04413_ _04678_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10991_ _00583_ clknet_leaf_40_clock net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08347__C _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08806__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09459__B _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10419__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _00017_ clknet_leaf_54_clock mem.mem_dff.code_mem\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06045__A1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10356_ _01793_ _05154_ _05157_ stack\[17\]\[1\] _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09782__A2 _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10569__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _04994_ _05093_ _05101_ stack\[30\]\[7\] _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08589__I _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09298__A1 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06837__I mem.mem_dff.code_mem\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05403__S0 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05400_ _00951_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06380_ _01890_ _01808_ _01916_ _01904_ _01917_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05331_ _00883_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08050_ _03253_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05262_ _00799_ _00814_ _00816_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07001_ _02371_ _02429_ _02425_ _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A1 _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__B1 _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__B2 stack\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06036__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_92_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__B1 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _03853_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07903_ _03136_ _03133_ _03137_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08883_ net151 _03948_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06013__S _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07834_ _02968_ _03074_ _03082_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05547__B1 stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07765_ _03027_ _03020_ _03029_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06716_ _02205_ _02202_ _02206_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09504_ _03281_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07696_ mem.mem_dff.code_mem\[31\]\[5\] _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _01027_ _04368_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06647_ _02150_ _02140_ _02151_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09366_ _04339_ _04344_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08962__I _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06578_ mem.mem_dff.code_mem\[2\]\[0\] _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08317_ mem.mem_dff.data_mem\[2\]\[5\] _03327_ _03329_ mem.mem_dff.data_mem\[6\]\[5\]
+ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05529_ _01043_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09297_ _04270_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08248_ mem.mem_dff.code_mem\[11\]\[3\] _03299_ _02443_ mem.mem_dff.code_mem\[13\]\[3\]
+ mem.mem_dff.code_mem\[26\]\[3\] _03300_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10711__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ mem.mem_dff.code_mem\[0\]\[1\] _03290_ _03373_ _03316_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09213__A1 stack\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10210_ _03868_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11190_ net235 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07775__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10374__A3 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ _04986_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput180 net180 o_wb_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_4_0_0_clock clknet_3_0_0_clock clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xoutput191 net191 rambus_wb_addr_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10072_ _01197_ _04935_ _04939_ net128 _04139_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10974_ _00566_ clknet_leaf_42_clock net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06266__A1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05510__B _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06392__I _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10062__A2 _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05313__I0 stack\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_114_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06018__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _00000_ clknet_leaf_139_clock stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06018__B2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _05061_ _05141_ _05146_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05736__I _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09208__I _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A2 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08715__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05880_ _00852_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07951__I _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09371__C _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _02847_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06501_ _01999_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ mem.mem_dff.code_mem\[25\]\[6\] _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10089__I _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _04169_ _04217_ _04219_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06432_ _01379_ _01397_ _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09151_ _03918_ _04166_ _04162_ _04167_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_188_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10734__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06363_ _01842_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08246__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09443__A1 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07398__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08102_ mem.mem_dff.code_mem\[9\]\[0\] _02321_ _02876_ mem.mem_dff.code_mem\[28\]\[0\]
+ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05314_ _00855_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05304__I0 stack\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ _03672_ _03993_ _01929_ _03192_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__09994__A2 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06008__S _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06294_ _01462_ _01482_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _03238_ _03210_ _03225_ stack\[28\]\[6\] _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05245_ _00769_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05855__I1 stack\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput60 i_wb_data[3] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput71 io_in[2] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput82 rambus_wb_dat_i[13] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput93 rambus_wb_dat_i[23] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10884__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08549__A3 _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__B1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09984_ _04866_ _01738_ _04868_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05646__I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09118__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05232__A2 _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _04006_ _04001_ _03999_ stack\[13\]\[2\] _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06980__A2 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08957__I _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08866_ _01796_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input21_I i_wb_addr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _02381_ _02135_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _03835_ _03899_ _03896_ stack\[6\]\[1\] _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _03015_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06477__I _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05381__I _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ mem.mem_dff.code_mem\[31\]\[1\] _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08485__A2 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__I _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06496__A1 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04388_ _04392_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _00282_ clknet_leaf_61_clock mem.mem_dff.data_mem\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ net91 _04291_ _04292_ net82 _04306_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__09434__A1 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06248__A1 _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06248__B2 _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__B1 _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05757__S _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09737__A2 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08945__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05556__I _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10124_ _04417_ _04961_ _04986_ _04592_ _04140_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10055_ net31 net30 net33 net32 _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10607__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08867__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09370__B1 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__I1 stack\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07920__A1 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_40_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05931__B1 _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10957_ _00549_ clknet_leaf_187_clock stack\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08476__A2 _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07720__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10283__A2 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10888_ _00480_ clknet_leaf_148_clock stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10035__A2 _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06239__B2 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09976__A2 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05837__I1 stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__I _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__B1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07739__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06411__B2 _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06981_ _02416_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05932_ _01302_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08720_ _03220_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09361__B1 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ _01796_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06014__I1 stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05863_ _01355_ _01400_ _01406_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07602_ _02901_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05415__B _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08582_ _03725_ _03730_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05794_ _01299_ _01336_ _01337_ _01304_ _01307_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_183_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07533_ _02847_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07464_ _02737_ _02792_ _02784_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10274__A2 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09401__I _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09203_ _01990_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06415_ _01937_ _01784_ _01951_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07395_ _02739_ _02733_ _02740_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _04129_ _04146_ _04153_ stack\[18\]\[4\] _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06346_ _01215_ _01737_ _01754_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08017__I _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07978__A1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _03758_ _04085_ _04093_ _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05828__I1 stack\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ _01814_ _01815_ _01816_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08016_ _03223_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input69_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06760__I mem.mem_dff.code_mem\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05228_ _00782_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05376__I _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _02004_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08918_ _03989_ _03991_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_131_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _04640_ _04645_ _04806_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output225_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _03770_ _03771_ _03197_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07902__A1 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ _00403_ clknet_leaf_171_clock stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10742_ _00334_ clknet_leaf_163_clock stack\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _00265_ clknet_leaf_60_clock mem.mem_dff.code_mem\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10017__A2 _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07969__A1 _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__A2 _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06641__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06670__I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09981__I _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11156_ _00748_ clknet_leaf_133_clock stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06944__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _04927_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11087_ _00679_ clknet_leaf_44_clock net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10038_ delay_counter\[6\] _04674_ _04899_ _01123_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07006__I mem.mem_dff.code_mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05950__S _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0_0_clock_I clknet_2_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09221__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06200_ _01736_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07180_ _02512_ _02565_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06880__A1 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06131_ _01652_ _01673_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07676__I _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06062_ _01603_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ net232 _02033_ _04481_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08924__A3 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__A1 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06935__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _04336_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05294__S1 _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06964_ _02401_ _02398_ _02402_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08137__A1 _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ _03820_ _03824_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06021__S _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05915_ stack\[30\]\[3\] stack\[31\]\[3\] _00821_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06895_ _02346_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09683_ delay_cycles\[23\] _04498_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09885__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09885__B2 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05846_ _01266_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08634_ _01588_ _03770_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_leaf_5_clock clknet_4_2_0_clock clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_215_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05860__S _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05777_ _00851_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08565_ _01827_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05910__A3 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ _02055_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__A2 _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08496_ _01893_ _03631_ _03660_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07447_ _02752_ _02776_ _02772_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06871__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ _02726_ _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09117_ _01638_ _03643_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06329_ _00839_ _01761_ _00916_ _00980_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08612__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10452__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06490__I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09048_ _04089_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output175_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _00602_ clknet_leaf_45_clock mem.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06926__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05985__I0 stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__B1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08679__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05362__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09628__B2 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05901__A3 _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06665__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10187__I _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10725_ _00317_ clknet_leaf_50_clock mem.mem_dff.data_mem\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05502__C _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06862__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10656_ _00248_ clknet_leaf_95_clock mem.mem_dff.code_mem\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ _00179_ clknet_leaf_81_clock mem.mem_dff.code_mem\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10136__B _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__S _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11139_ _00731_ clknet_leaf_193_clock stack\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08120__I _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09867__A1 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09867__B2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05700_ _01241_ _01243_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06680_ _02144_ _02176_ _02166_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05631_ _01171_ _01172_ _01177_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08350_ _03539_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10229__A2 _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05562_ _01102_ _01107_ _01110_ _01053_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07301_ _02666_ _02663_ _02667_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08281_ _02015_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05493_ _01015_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08842__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10475__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _02127_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_4_0_clock_I clknet_3_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _02556_ _02549_ _02559_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06114_ _01654_ _01655_ _01656_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05259__I2 stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10401__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07094_ _02036_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06016__S _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_162_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06045_ _01574_ _01231_ _01102_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout236 net217 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ net153 _04740_ _04741_ _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xfanout247 net248 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout258 net159 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11100__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _03207_ _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09735_ cycles_per_ms\[23\] cycles_per_ms\[22\] cycles_per_ms\[21\] cycles_per_ms\[20\]
+ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06947_ _02389_ _02386_ _02378_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_153_clock clknet_4_5_0_clock clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09666_ delay_cycles\[20\] _04496_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06878_ _02322_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08530__A1 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08530__B2 stack\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08617_ _03757_ _03759_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05344__A1 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05829_ _01363_ _01370_ _01372_ _00803_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09597_ _04556_ _04490_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_87_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06485__I _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10818__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08548_ _03191_ _03639_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_165_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_168_clock clknet_4_3_0_clock clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _03633_ _03642_ _03648_ stack\[19\]\[0\] _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__A1 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10510_ _00102_ clknet_leaf_110_clock mem.mem_dff.code_mem\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__C _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _00033_ clknet_leaf_67_clock mem.mem_dff.code_mem\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10968__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10372_ _03858_ _03188_ _03189_ _03702_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06072__A2 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05765__S _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_106_clock clknet_4_13_0_clock clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__S _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10156__A1 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09010__A2 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05564__I _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09849__A1 _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08521__A1 _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10498__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__B1 _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06835__A1 _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _00300_ clknet_leaf_37_clock mem.mem_dff.data_mem\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10639_ _00231_ clknet_leaf_103_clock mem.mem_dff.code_mem\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08588__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10395__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11123__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__A2 _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10147__A1 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05249__S1 _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _03065_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_70_clock clknet_4_14_0_clock clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08760__A1 stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06801_ _02259_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07781_ mem.mem_dff.data_mem\[2\]\[0\] _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 i_la_addr[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09520_ _04477_ _04480_ _04402_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06732_ mem.mem_dff.code_mem\[5\]\[6\] _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09390__B _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_109_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09451_ _04418_ _04384_ _04421_ _04422_ _04401_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06663_ net233 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10967__D _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_85_clock clknet_4_15_0_clock clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_213_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08402_ net123 _03112_ _03578_ _03579_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05614_ _01103_ _01161_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05421__S1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05423__B _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05877__A2 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09382_ net128 _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06594_ net244 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09068__A2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08333_ _03517_ _03520_ _03521_ _03522_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05545_ _00934_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ _03452_ _03453_ _03454_ _03455_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06826__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05476_ _01026_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07215_ _02557_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08195_ _02926_ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07146_ _02512_ _02539_ _02546_ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10386__A1 _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23_clock clknet_4_10_0_clock clknet_leaf_23_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07077_ mem.mem_dff.code_mem\[14\]\[6\] _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07864__I _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input51_I i_wb_data[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01528_ _01542_ _01556_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_clock clknet_4_9_0_clock clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspell_261 o_wb_data[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output138_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07979_ _01710_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09718_ _04677_ _01244_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10640__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _00582_ clknet_leaf_41_clock mem.select vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08503__A1 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _04578_ _04607_ _04608_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09059__A2 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08267__B1 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10790__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06117__I0 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08363__C _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07490__A1 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11146__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10424_ _00016_ clknet_leaf_54_clock mem.mem_dff.code_mem\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A1 _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06045__A2 _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10355_ _03890_ _05152_ _05158_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10129__A1 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10286_ _03908_ _05105_ _05106_ _05107_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10129__B2 _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_215_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09534__A3 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07723__B _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_110_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10301__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05403__S1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07014__I _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05330_ _00767_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06853__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__C _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05261_ _00815_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10375__I _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07000_ mem.mem_dff.code_mem\[12\]\[5\] _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_200_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__A1 _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10368__B2 stack\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06036__A2 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _03846_ _04017_ _04018_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08981__B2 stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07902_ _03107_ _03134_ _03127_ _03137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08882_ stack\[26\]\[6\] _03950_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07833_ _03065_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05547__A1 _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05547__B2 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07764_ _02968_ _03021_ _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09404__I _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09503_ _00850_ _04449_ _04466_ _04467_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06715_ _02144_ _02203_ _02195_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07695_ _02971_ _02972_ _02974_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04406_ _04404_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06646_ _02129_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09365_ mem.io_data_out\[6\] _04267_ _04343_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06577_ _02091_ _02084_ _02093_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_209_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ mem.mem_dff.data_mem\[4\]\[5\] _03323_ _03324_ mem.mem_dff.data_mem\[5\]\[5\]
+ _03325_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_162_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input99_I rambus_wb_dat_i[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05528_ _01042_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09296_ _03099_ _04279_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__A3 _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _03436_ _03437_ _03438_ _03439_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05459_ _00767_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05600__C _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08178_ _03338_ _03339_ _03348_ _03372_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_134_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10359__A1 _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09213__A2 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06027__A2 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ net187 _02023_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ net183 _04999_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08972__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput170 net170 o_wb_data[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput181 net181 o_wb_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput192 net192 rambus_wb_clk_o vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_121_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10071_ _04938_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08185__C1 mem.mem_dff.data_mem\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__C _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10973_ _00565_ clknet_leaf_43_clock net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06673__I _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05313__I1 stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05289__I _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ _03854_ _05193_ _05195_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10338_ _01888_ _05132_ _05145_ stack\[16\]\[4\] _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A3 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10269_ _05091_ _05096_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08715__A1 _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09224__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09140__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06500_ _02028_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07480_ _02805_ _02802_ _02806_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _01949_ _01940_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05701__A1 _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07679__I mem.mem_dff.code_mem\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ _00842_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06362_ _01772_ _01899_ _01890_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09443__A2 _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03291_ _03294_ _03295_ _03296_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05313_ stack\[15\]\[1\] stack\[12\]\[1\] stack\[13\]\[1\] stack\[14\]\[1\] _00857_
+ _00847_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09081_ _04114_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06293_ _01722_ net60 _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_30_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05304__I1 stack\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05465__B1 stack\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05244_ _00798_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08032_ _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 i_wb_data[16] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05855__I2 stack\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput61 i_wb_data[4] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput72 io_in[3] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput83 rambus_wb_dat_i[14] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10980__D _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput94 rambus_wb_dat_i[24] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_192_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08549__A4 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08954__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__B2 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__S _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _02031_ _04867_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08934_ _01824_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08167__C1 mem.mem_dff.code_mem\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ _03952_ _03943_ _03953_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07816_ mem.mem_dff.data_mem\[3\]\[0\] _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10409__CLK clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08796_ _03891_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06193__A1 _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input14_I i_la_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07747_ _02381_ _03014_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05940__A1 _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__B1 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ _02955_ _02959_ _02961_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09682__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10559__CLK clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09417_ _00919_ _04368_ _04389_ _04391_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06629_ _02136_ _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06496__A2 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ net105 _04304_ _02134_ net99 _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _04263_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09198__B2 stack\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09737__A3 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06442__B _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08945__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08945__B2 stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10123_ _04949_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10054_ net35 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09370__A1 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07273__B _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__B2 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07920__A2 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05931__A1 _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_0_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05931__B2 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10268__B1 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _00548_ clknet_leaf_187_clock stack\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10887_ _00479_ clknet_leaf_143_clock stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__S0 _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07436__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05948__S _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09189__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__B2 stack\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05747__I _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07739__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08936__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08123__I _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06411__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06980_ _02411_ _02415_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07962__I _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I i_la_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _00794_ _01473_ _01474_ _01363_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A1 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09361__B2 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ _03785_ _03775_ _03786_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05862_ _01401_ _01402_ _01404_ _01405_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _02787_ _02440_ _02198_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__C _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ stack\[31\]\[5\] _03727_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05793_ stack\[20\]\[0\] stack\[21\]\[0\] _00811_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05922__A1 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09113__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05922__B2 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__B1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07532_ _02847_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08793__I _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09664__A2 _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ mem.mem_dff.code_mem\[25\]\[1\] _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06478__A2 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09202_ _04133_ _04203_ _04204_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06414_ _01122_ _01785_ _01949_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10851__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07394_ _02710_ _02734_ _02727_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09133_ _04056_ _04144_ _04154_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06345_ _01801_ _01876_ _01880_ _01883_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05858__S _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07978__A2 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09064_ _00983_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06276_ exec.memory_input\[2\] _01744_ _01779_ _00877_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_191_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05989__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05989__B2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05227_ _00774_ _00775_ _00768_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_08015_ _01886_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09966_ _04850_ _04856_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05610__B1 stack\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08848_ _03936_ _03934_ _03938_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output120_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05913__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ _03846_ _03885_ _03886_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output218_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05913__B2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_157_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _00402_ clknet_leaf_166_clock stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__C1 mem.mem_dff.code_mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10741_ _00333_ clknet_leaf_134_clock stack\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10672_ _00264_ clknet_leaf_60_clock mem.mem_dff.code_mem\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09748__B intr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09467__C _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ _00747_ clknet_leaf_190_clock stack\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09483__B _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10106_ _01228_ _04969_ _04941_ _04281_ _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_11086_ _00678_ clknet_leaf_10_clock net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10724__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10037_ _04903_ _04904_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05904__A1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10874__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09646__A2 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09502__I _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07657__A1 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10939_ _00531_ clknet_leaf_183_clock stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_4_0_clock_I clknet_2_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ _00850_ _01671_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08082__A1 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06061_ _01598_ _01604_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05477__I _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08909__A1 stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09820_ _04752_ _04744_ _04754_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__I _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09751_ intr_enable\[0\] _04706_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06963_ _02371_ _02399_ _02395_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05994__I1 stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08702_ _03823_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05914_ stack\[28\]\[3\] stack\[29\]\[3\] _01417_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09682_ _04250_ _04641_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06894_ _02345_ _02319_ _02096_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09885__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08633_ _01616_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05845_ _01259_ _01388_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08564_ stack\[31\]\[3\] _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05371__A2 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05776_ _01297_ _01308_ _01314_ _01319_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09412__I _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07515_ mem.mem_dff.code_mem\[26\]\[5\] _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08495_ _03659_ _03641_ _03657_ stack\[19\]\[5\] _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ mem.mem_dff.code_mem\[24\]\[6\] _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07377_ _02613_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input81_I rambus_wb_dat_i[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09116_ _03282_ _04141_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10404__B1 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06328_ _01842_ _01772_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_202_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _03740_ _04085_ _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06259_ _01722_ net59 _01799_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10747__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08698__I _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09949_ _04840_ _04845_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05985__I1 stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__A1 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__B2 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06139__A1 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06946__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09628__A2 _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _00316_ clknet_leaf_51_clock mem.mem_dff.data_mem\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10655_ _00247_ clknet_leaf_95_clock mem.mem_dff.code_mem\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08064__A1 mem.io_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10586_ _00178_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__B1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06378__A1 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10174__A2 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_clock_I clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11138_ _00730_ clknet_leaf_187_clock stack\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08119__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11069_ _00661_ clknet_opt_1_0_clock net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09867__A2 _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07878__A1 _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05630_ net189 net188 _01176_ net190 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_184_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05760__I _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11052__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05561_ _01103_ _01108_ _01109_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10378__I _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07300_ _02608_ _02664_ _02660_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08280_ _03461_ _03469_ _03470_ _03471_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_05492_ _01012_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07231_ mem.mem_dff.code_mem\[18\]\[7\] _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_203_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07687__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07162_ _02527_ _02550_ _02558_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08055__A1 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08055__B2 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_105_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06113_ net1 net2 net17 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07093_ mem.mem_dff.code_mem\[15\]\[1\] _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_4_8_0_clock_I clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05259__I3 stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06044_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__A2 _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout237 net239 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_09803_ _01827_ _04732_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07030__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout248 net211 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07995_ _01756_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09307__A1 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ cycles_per_ms\[19\] _04517_ _04514_ cycles_per_ms\[16\] _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09307__B2 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06946_ _02143_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09665_ cycles_per_ms\[20\] _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06877_ mem.mem_dff.code_mem\[9\]\[4\] _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07371__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__A2 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08616_ _03758_ _03742_ _03749_ net147 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05828_ stack\[26\]\[7\] stack\[27\]\[7\] _01371_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ delay_cycles\[7\] _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05344__A2 _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08547_ _01683_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05759_ _01302_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08478_ _03647_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08294__B2 mem.mem_dff.code_mem\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _02737_ _02765_ _02756_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06844__A2 _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07597__I _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _00032_ clknet_leaf_68_clock mem.mem_dff.code_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__A1 _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10371_ _04137_ _05165_ _05151_ _03855_ _05167_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_136_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__B2 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__A2 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09849__A2 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11075__CLK clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09480__C _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06676__I _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08891__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08285__B2 mem.mem_dff.data_mem\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05718__S0 _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10092__A1 _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _00299_ clknet_leaf_30_clock mem.mem_dff.data_mem\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08037__A1 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10638_ _00230_ clknet_leaf_103_clock mem.mem_dff.code_mem\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06117__S _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ _00161_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10395__A2 _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05755__I _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08131__I _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06800_ mem.mem_dff.code_mem\[7\]\[4\] _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ _03038_ _03031_ _03040_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06771__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07970__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 i_la_addr[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_06731_ _02216_ _02213_ _02217_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08512__A2 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09450_ _04334_ _04399_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06662_ mem.mem_dff.code_mem\[3\]\[7\] _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10442__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06586__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05490__I _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ net123 _03573_ _03576_ _03112_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05613_ _01077_ stack\[24\]\[7\] stack\[25\]\[7\] _01150_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _01222_ _04315_ _04358_ _04337_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06593_ mem.mem_dff.code_mem\[2\]\[2\] _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09897__I _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08332_ mem.mem_dff.code_mem\[7\]\[6\] _03428_ _02443_ mem.mem_dff.code_mem\[13\]\[6\]
+ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05544_ _00932_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10592__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ mem.mem_dff.code_mem\[6\]\[4\] _02226_ _02927_ mem.mem_dff.code_mem\[30\]\[4\]
+ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05475_ _01025_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07214_ mem.mem_dff.code_mem\[18\]\[3\] _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _02225_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07145_ _02494_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10386__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07076_ _02488_ _02484_ _02490_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05262__A1 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06027_ _01563_ _01570_ _01357_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I i_wb_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__A1 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11098__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _01699_ _01703_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xspell_262 o_wb_data[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09717_ single_step _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06929_ _02373_ _02364_ _02374_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09700__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ _04572_ _04573_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__A2 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output200_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ _04529_ _04531_ _04536_ _04538_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10935__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06117__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__A1 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07490__A2 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07120__I mem.mem_dff.code_mem\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10423_ _00015_ clknet_leaf_54_clock mem.mem_dff.code_mem\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10354_ _01758_ _05154_ _05157_ stack\[17\]\[0\] _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05253__A1 _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10285_ _03238_ _05093_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10129__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05575__I _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05508__C _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08742__A2 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10465__CLK clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10301__A2 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05939__S0 _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05867__I0 stack\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05260_ _00773_ _00782_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_179_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09758__A1 _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_152_clock clknet_4_5_0_clock clknet_leaf_152_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06036__A3 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08430__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08950_ _03851_ _03997_ _04009_ stack\[13\]\[6\] _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08981__A2 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__CLK clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ mem.mem_dff.data_mem\[5\]\[1\] _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08881_ _01933_ _03964_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_167_clock clknet_4_3_0_clock clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07832_ mem.mem_dff.data_mem\[3\]\[3\] _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07914__B _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05547__A2 stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07763_ _03010_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10978__D _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10958__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09502_ _04336_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06714_ mem.mem_dff.code_mem\[5\]\[1\] _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07694_ _02943_ _02973_ _02969_ _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09694__B1 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ net154 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06645_ _02149_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08249__A1 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09364_ _04340_ _04341_ _04342_ _04274_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06576_ _02064_ _02085_ _02092_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_105_clock clknet_4_13_0_clock clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08315_ mem.mem_dff.data_mem\[1\]\[5\] _03016_ _03070_ mem.mem_dff.data_mem\[3\]\[5\]
+ mem.mem_dff.data_mem\[7\]\[5\] _03321_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_127_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05527_ _00960_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09295_ net95 net230 net229 net86 net228 net109 _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_178_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05858__I0 stack\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08246_ mem.mem_dff.code_mem\[17\]\[3\] _02562_ _02620_ mem.mem_dff.code_mem\[19\]\[3\]
+ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05458_ _00924_ _00959_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09749__A1 _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08177_ _03361_ _03371_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05389_ _00940_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10359__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07128_ _02531_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07096__B _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ mem.mem_dff.code_mem\[14\]\[2\] _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08972__A2 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10007__S _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput160 net160 o_wb_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10488__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput171 net171 o_wb_data[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput182 net182 o_wb_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput193 net193 rambus_wb_cyc_o vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10070_ _04936_ _04937_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10972_ _00564_ clknet_4_3_0_clock net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08488__A1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08488__B2 stack\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11113__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_6_0_clock clknet_4_12_0_clock clknet_opt_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09330__I _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09988__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__I0 stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__B1 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05313__I2 stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10406_ _04994_ _05188_ _05191_ stack\[15\]\[7\] _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08412__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08412__B2 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_84_clock clknet_4_15_0_clock clknet_leaf_84_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08963__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10337_ _05134_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10268_ _04915_ _05093_ _05095_ stack\[30\]\[0\] _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08715__A2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10199_ _04483_ _04956_ _05037_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_clock clknet_4_13_0_clock clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08479__A1 _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__B2 stack\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09140__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10286__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_22_clock clknet_4_10_0_clock clknet_leaf_22_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07151__A1 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _01934_ _01964_ _01965_ _01966_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06864__I _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09240__I _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A1 _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__B2 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _01025_ _01868_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08100__B1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08100_ mem.mem_dff.code_mem\[6\]\[0\] _02226_ _02927_ mem.mem_dff.code_mem\[30\]\[0\]
+ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_37_clock clknet_4_11_0_clock clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05312_ _00819_ _00865_ _00807_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09080_ _03820_ _03941_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06292_ _01767_ _01831_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05304__I2 stack\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05465__A1 _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08031_ _01123_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput40 i_wb_addr[8] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_05243_ _00783_ _00797_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05465__B2 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07909__B _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput51 i_wb_data[17] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05855__I3 stack\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput62 i_wb_data[5] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__10630__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput73 io_in[4] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07206__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput84 rambus_wb_dat_i[15] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_196_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 rambus_wb_dat_i[25] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08954__A2 _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09982_ _04865_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _03952_ _04003_ _04005_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06104__I _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ _03835_ _03947_ _03950_ stack\[26\]\[1\] _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07815_ _03064_ _03057_ _03067_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _03890_ _03892_ _03897_ _03900_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05240__I1 stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07746_ _00762_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11136__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05940__A2 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07677_ _02930_ _02960_ _02953_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07142__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09416_ _04386_ _04390_ _04367_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06628_ _02133_ _02135_ _02095_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06774__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09150__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09347_ _01186_ _04315_ _04327_ _04289_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06559_ mem.mem_dff.code_mem\[1\]\[3\] _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _03621_ _04255_ _04262_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_201_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output198_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08229_ mem.mem_dff.code_mem\[23\]\[3\] _03391_ _03392_ mem.mem_dff.code_mem\[31\]\[3\]
+ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_0_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09198__A2 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_153_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09737__A4 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06442__C _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__A2 _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10122_ _04984_ _04985_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09753__C _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06008__I0 stack\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10053_ net36 _04916_ _04920_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06949__I mem.mem_dff.code_mem\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09370__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06184__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A1 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10503__CLK clknet_leaf_107_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _00547_ clknet_leaf_183_clock stack\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07133__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _00478_ clknet_leaf_146_clock stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08881__A1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09060__I _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05790__S1 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10653__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05447__A1 _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05998__A2 _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09189__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08404__I _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08936__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06947__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05930_ stack\[0\]\[3\] stack\[1\]\[3\] _01438_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11159__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05763__I _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09361__A2 _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05861_ _01271_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ mem.mem_dff.code_mem\[29\]\[0\] _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _03728_ _03700_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05792_ stack\[22\]\[0\] stack\[23\]\[0\] _00882_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05383__B1 _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10259__A1 _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07531_ _02759_ _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09113__A2 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10259__B2 stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07124__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ _02786_ _02791_ _02793_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09201_ _04135_ _04193_ _04200_ stack\[20\]\[6\] _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06413_ _01123_ _01949_ _01735_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07393_ mem.mem_dff.code_mem\[23\]\[2\] _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09132_ _04126_ _04147_ _04153_ stack\[18\]\[3\] _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06344_ _01743_ _01881_ _01882_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05438__A1 _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ stack\[23\]\[3\] _04090_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06275_ _01736_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ _01829_ _03213_ _03222_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05226_ _00780_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05874__S _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09965_ _04485_ _04854_ _04852_ _04508_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05610__A1 _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05610__B2 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07374__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08916_ _01605_ _03771_ _03821_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09896_ _04338_ _04803_ _04804_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05673__I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08189__C _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _03937_ _03930_ _03928_ stack\[7\]\[7\] _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _03851_ _03865_ _03872_ stack\[11\]\[6\] _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09104__A2 _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output113_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07729_ _02116_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08312__B1 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__C2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10676__CLK clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _00332_ clknet_leaf_160_clock stack\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10671_ _00263_ clknet_leaf_59_clock mem.mem_dff.code_mem\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08918__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09040__A1 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _00746_ clknet_leaf_191_clock stack\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10105_ _04956_ _04970_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11085_ _00677_ clknet_leaf_10_clock net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05583__I _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10036_ _04884_ _04905_ _04906_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05516__C _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05904__A2 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08303__B1 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10938_ _00530_ clknet_leaf_180_clock stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10869_ _00461_ clknet_leaf_140_clock stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08606__A1 stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07973__I _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05279__S0 _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10549__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06962_ mem.mem_dff.code_mem\[11\]\[5\] _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09750_ _03618_ _04361_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05493__I _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08701_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05913_ _01409_ _01455_ _01456_ _01414_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09681_ net142 _04252_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06893_ _02287_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08542__B1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _01598_ _01604_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05844_ stack\[2\]\[7\] stack\[3\]\[7\] stack\[0\]\[7\] stack\[1\]\[7\] _00856_ _00869_
+ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07896__A2 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_101_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08563_ _01315_ _03706_ _03714_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05775_ _01299_ _01317_ _01318_ _01304_ _01279_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ _02829_ _02830_ _02833_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input109_I rambus_wb_dat_i[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _03227_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07445_ _02778_ _02775_ _02779_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05869__S _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ mem.mem_dff.code_mem\[22\]\[7\] _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _04140_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10404__A1 _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06327_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10404__B2 stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05668__I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input74_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09046_ _03743_ _04087_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08044__I _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06258_ _01724_ _01798_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05209_ _00763_ _00764_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09022__A1 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06189_ _01230_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06387__A2 _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06499__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09948_ _04532_ _04835_ _04843_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05985__I2 stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__A2 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output230_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09879_ _04791_ _04793_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__B1 _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10723_ _00315_ clknet_leaf_50_clock mem.mem_dff.data_mem\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06311__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05779__S _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10654_ _00246_ clknet_leaf_94_clock mem.mem_dff.code_mem\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10585_ _00177_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09261__B2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05578__I _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09013__A1 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07793__I mem.mem_dff.data_mem\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07575__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06378__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ _00729_ clknet_leaf_184_clock stack\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10841__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A3 _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11068_ _00660_ clknet_4_0_0_clock net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ delay_counter\[2\] _04888_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_4_15_0_clock_I clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07878__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10331__B1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10991__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05560_ _01093_ stack\[27\]\[6\] _01094_ stack\[26\]\[6\] _01051_ _01109_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08129__I _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05491_ _01009_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07230_ _02610_ _02603_ _02611_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _02557_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10394__I stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06112_ net18 net29 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06066__A1 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07092_ _02497_ _02501_ _02503_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ _01254_ _01257_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07917__B _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09555__A2 _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09802_ _04723_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout238 net239 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07994_ stack\[28\]\[0\] _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout249 net250 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06945_ mem.mem_dff.code_mem\[11\]\[1\] _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09733_ _01189_ _01194_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09664_ _04528_ _04620_ _04622_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_06876_ _02330_ _02323_ _02332_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05424__S0 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05827_ _00855_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08615_ _03220_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09595_ delay_cycles\[8\] _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05758_ _01265_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08546_ _03699_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ _03185_ _03641_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09491__A1 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05689_ _01184_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ mem.mem_dff.code_mem\[24\]\[1\] _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06782__I _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09298__C _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10714__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__B _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07359_ mem.mem_dff.code_mem\[22\]\[3\] _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05398__I _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06057__A1 _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output180_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10370_ stack\[17\]\[7\] _05157_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09029_ _04006_ _04070_ _04074_ stack\[9\]\[2\] _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05804__A1 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__B1 _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08285__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__S1 _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06296__A1 _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10706_ _00298_ clknet_leaf_29_clock mem.mem_dff.data_mem\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10637_ _00229_ clknet_leaf_102_clock mem.mem_dff.code_mem\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08037__A2 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09234__A1 _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__A1 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10568_ _00160_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09785__A2 _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10499_ _00091_ clknet_leaf_108_clock mem.mem_dff.code_mem\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05559__B1 stack\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05972__S _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06730_ _02122_ _02214_ _02210_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 i_la_addr[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10304__B1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05771__I stack\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__I _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08287__C _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06661_ _02159_ _02154_ _02162_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10389__I stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08400_ _03581_ _03584_ _03585_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_149_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05612_ _01141_ _01158_ _01159_ _01134_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _04303_ _04353_ _04357_ _04263_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06592_ _02105_ _02100_ _02106_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08331_ mem.mem_dff.code_mem\[9\]\[6\] _02320_ _02468_ mem.mem_dff.code_mem\[14\]\[6\]
+ mem.mem_dff.code_mem\[28\]\[6\] _03430_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05543_ _01041_ _01091_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_205_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08262_ mem.mem_dff.code_mem\[15\]\[4\] _02499_ _02902_ mem.mem_dff.code_mem\[29\]\[4\]
+ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05474_ _01024_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07213_ _02596_ _02590_ _02598_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05885__I1 stack\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ mem.mem_dff.code_mem\[15\]\[2\] _02499_ _02902_ mem.mem_dff.code_mem\[29\]\[2\]
+ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07144_ mem.mem_dff.code_mem\[16\]\[3\] _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10887__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09846__C _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07647__B _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07075_ _02489_ _02486_ _02481_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06551__B _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06026_ _01282_ _01566_ _01569_ _01307_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_195_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08736__B1 _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input37_I i_wb_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ _01691_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xspell_263 o_wb_data[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09716_ _04412_ _01240_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06928_ _02279_ _02367_ _02361_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09153__I _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__A2 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _04581_ _04595_ _04602_ _04605_ _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _02318_ _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07711__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05317__A3 _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _04537_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_208_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08529_ _03681_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08267__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09464__A1 _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06278__A1 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10074__A2 _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07401__I mem.mem_dff.code_mem\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08019__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11070__D _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__A1 _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__A3 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10422_ _00014_ clknet_leaf_53_clock mem.mem_dff.code_mem\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _05156_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05253__A2 _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10284_ stack\[30\]\[6\] _05095_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11042__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_2_0_clock clknet_4_2_0_clock clknet_opt_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05792__S _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__A1 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05939__S1 _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_148_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A1 _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A1 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05316__I0 stack\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08407__I _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05867__I1 stack\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09758__A2 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07769__A1 _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06441__A1 _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__B1 _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07900_ _03129_ _03133_ _03135_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08880_ _01931_ _03231_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07831_ _03078_ _03072_ _03080_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07941__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07762_ mem.mem_dff.data_mem\[1\]\[3\] _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _04382_ _01588_ _04438_ _04465_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06713_ _02197_ _02202_ _02204_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07693_ _02958_ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09694__A1 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09694__B2 _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09432_ net154 _04404_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06644_ net242 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06575_ _02065_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09363_ _01172_ mem.dff_data_out\[6\] _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08314_ mem.mem_dff.code_mem\[0\]\[5\] _03451_ _03495_ _03504_ _03473_ _03505_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10056__A2 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05526_ _01075_ net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_178_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09294_ _01212_ _04265_ _04278_ _03627_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09997__A2 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ mem.mem_dff.code_mem\[1\]\[3\] _02071_ _03405_ mem.mem_dff.code_mem\[16\]\[3\]
+ _02027_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05858__I1 stack\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05457_ _00972_ _01003_ _01007_ _00974_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06680__A1 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08176_ _03362_ _03363_ _03367_ _03370_ _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09749__A2 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05388_ _00790_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _02016_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08421__A2 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06432__A1 _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07058_ _02475_ _02471_ _02476_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput150 net150 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput161 net161 o_wb_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_161_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06983__A2 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput172 net172 o_wb_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06009_ stack\[28\]\[1\] stack\[29\]\[1\] _01438_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput183 net183 o_wb_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput194 net194 rambus_wb_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08185__A1 mem.mem_dff.data_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08185__B2 mem.mem_dff.data_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07932__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10902__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__B1 _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10971_ _00563_ clknet_leaf_43_clock net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08488__A2 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07840__B _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_clock clknet_4_0_0_clock clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09437__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05360__B _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A1 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__B2 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__I1 stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05313__I3 stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05787__S _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06970__I _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10405_ _03963_ _05193_ _05194_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10432__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05586__I _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08963__A3 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10336_ _05059_ _05141_ _05144_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_74_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09912__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10582__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10198_ net176 _05035_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07306__I _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__B1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__A2 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09676__B2 _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__A4 delay_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10038__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ _01873_ _01897_ _01874_ _01871_ _01866_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11088__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05311_ stack\[7\]\[1\] stack\[4\]\[1\] stack\[5\]\[1\] stack\[6\]\[1\] _00832_ _00823_
+ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06291_ net11 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05304__I3 stack\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07976__I _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08030_ _03232_ _03235_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05242_ _00787_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05465__A2 stack\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 i_wb_addr[20] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09396__C _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput41 i_wb_addr[9] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput52 i_wb_data[18] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 i_wb_data[6] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08939__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput74 io_in[5] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput85 rambus_wb_dat_i[16] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput96 rambus_wb_dat_i[26] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06414__A1 _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04865_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10925__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ _04004_ _04001_ _03999_ stack\[13\]\[1\] _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08167__A1 mem.mem_dff.code_mem\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__B2 mem.mem_dff.code_mem\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06017__I1 stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10989__D _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _01763_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A1 _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07814_ _02981_ _03058_ _03066_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08794_ _03898_ _03899_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05240__I2 stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ mem.mem_dff.data_mem\[1\]\[0\] _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10277__A2 _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ _02958_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09415_ net139 _04378_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06627_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06350__B1 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06558_ _02078_ _02073_ _02079_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09346_ _04303_ _04322_ _04326_ _04301_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05509_ stack\[7\]\[5\] stack\[4\]\[5\] stack\[5\]\[5\] stack\[6\]\[5\] _01029_ _00969_
+ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06489_ _02020_ net227 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09277_ _01661_ _04259_ _04261_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_194_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10455__CLK clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ mem.mem_dff.code_mem\[6\]\[3\] _03388_ _03389_ mem.mem_dff.code_mem\[30\]\[3\]
+ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ mem.mem_dff.code_mem\[5\]\[1\] _03352_ _03353_ mem.mem_dff.code_mem\[20\]\[1\]
+ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06956__A2 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ net179 _04957_ _04429_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__I1 stack\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10052_ net37 _04919_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07905__A1 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_151_clock clknet_4_5_0_clock clknet_leaf_151_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10268__A2 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ _00546_ clknet_leaf_179_clock stack\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__A1 mem.mem_dff.code_mem\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10885_ _00477_ clknet_leaf_143_clock stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08881__A2 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_166_clock clknet_4_3_0_clock clknet_leaf_166_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05447__A2 _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__A1 _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06205__I _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06947__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10319_ _04137_ _05129_ _05117_ _04112_ _05131_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_98_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_clock clknet_4_13_0_clock clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05860_ stack\[22\]\[6\] stack\[23\]\[6\] _01403_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07036__I mem.mem_dff.code_mem\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05980__S _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05791_ _01260_ _01334_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05383__A1 _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_119_clock clknet_4_12_0_clock clknet_leaf_119_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07530_ _02845_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ _02704_ _02792_ _02784_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10478__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ _03235_ _04109_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06412_ _01935_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06883__A1 _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07392_ _02736_ _02733_ _02738_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05930__I0 stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _04148_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06343_ _01074_ _01745_ _01780_ _00983_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__B1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08624__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09062_ _04099_ _04101_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06274_ _01746_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05225_ _00772_ _00777_ _00779_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08013_ _03221_ _03209_ _03205_ stack\[28\]\[3\] _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__A1 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09854__C _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09964_ _04850_ _04855_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11103__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ _03669_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05610__A2 stack\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09895_ _01624_ _01590_ _04648_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08846_ _01170_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08777_ _03664_ _03849_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05989_ _01390_ _01531_ _01532_ _01394_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07728_ _02998_ _02991_ _03000_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09161__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08312__B2 mem.mem_dff.code_mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07659_ mem.mem_dff.code_mem\[30\]\[5\] _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _00262_ clknet_leaf_59_clock mem.mem_dff.code_mem\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__I0 stack\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09329_ _04267_ _04309_ _04310_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09812__A1 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_clock clknet_4_13_0_clock clknet_leaf_98_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A2 _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_clock clknet_4_8_0_clock clknet_leaf_21_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06929__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _00745_ clknet_leaf_175_clock stack\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05864__I _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10104_ _04603_ _04963_ _04944_ _01133_ net257 _04939_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_11084_ _00676_ clknet_leaf_129_clock net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09879__A1 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10035_ delay_counter\[5\] _04882_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09780__B _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36_clock clknet_4_10_0_clock clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08551__A1 _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05904__A3 _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06909__B _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10620__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A1 mem.mem_dff.code_mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08303__B2 mem.mem_dff.code_mem\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _00529_ clknet_leaf_149_clock stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06865__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05912__I0 stack\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10868_ _00460_ clknet_leaf_190_clock stack\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10770__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09803__A1 _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__A2 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _00391_ clknet_leaf_134_clock stack\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11126__CLK clknet_leaf_158_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05975__S _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__A1 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05279__S1 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06961_ _02397_ _02398_ _02400_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _03770_ _03771_ _03821_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05912_ stack\[24\]\[3\] stack\[25\]\[3\] _01412_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09680_ _04484_ _04499_ _04506_ _04638_ _04639_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06892_ mem.mem_dff.code_mem\[10\]\[0\] _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08542__A1 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__B2 stack\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ _03736_ _03767_ _03769_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05356__A1 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05843_ _01380_ _01383_ _01386_ _01306_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _03218_ _03711_ _03713_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09098__A2 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05774_ stack\[28\]\[2\] stack\[29\]\[2\] _00882_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07513_ _02831_ _02832_ _02827_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08493_ _01861_ _03631_ _03658_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07444_ _02721_ _02776_ _02772_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07375_ _02723_ _02716_ _02724_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06554__B _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04139_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06326_ _01498_ _01513_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10404__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06084__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _04086_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06257_ net10 _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05208_ mem.mem_dff.memory_type_data _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05885__S _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I i_wb_stb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10168__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06188_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09022__A2 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A1 stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08060__I _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09947_ _04532_ _04546_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__05595__A1 _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05985__I3 stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08995__I _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _04517_ _04792_ _04788_ net52 _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10643__CLK clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output223_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08829_ _03755_ _03919_ _03920_ net146 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__A1 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__B2 stack\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10793__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11073__D _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _00314_ clknet_leaf_30_clock mem.mem_dff.data_mem\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06847__A1 _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10653_ _00245_ clknet_leaf_94_clock mem.mem_dff.code_mem\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11149__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08235__I _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _00176_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09261__A2 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06075__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09013__A2 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08772__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _00728_ clknet_leaf_179_clock stack\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08119__A4 _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11067_ _00659_ clknet_opt_2_0_clock net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10018_ _04890_ _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout254_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05490_ _00972_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05510__A1 _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__I _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ _02376_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08145__I _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10516__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06111_ net17 _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_173_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07091_ _02472_ _02502_ _02495_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09685__B _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06042_ _01126_ _01576_ _01580_ _01321_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09004__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10666__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout239 net215 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07993_ _03204_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _01624_ _01590_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__B _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ _02380_ _02385_ _02387_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09663_ _04524_ _04525_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06875_ _02269_ _02324_ _02331_ _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10322__A1 _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ stack\[3\]\[3\] _03746_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05826_ stack\[24\]\[7\] stack\[25\]\[7\] _01369_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05424__S1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09594_ cycles_per_ms\[8\] _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08279__B1 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08545_ _03194_ _03195_ _03197_ _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_05757_ stack\[20\]\[2\] stack\[21\]\[2\] _00901_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06829__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _03643_ _03645_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05688_ _01231_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _02758_ _02764_ _02766_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07358_ _02709_ _02703_ _02711_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06309_ _01816_ _01847_ _01848_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _02657_ _02652_ _02658_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _04050_ _04068_ _04076_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05804__A2 stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output173_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05568__A1 _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11068__D _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05568__B2 stack\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08506__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10313__A1 stack\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09482__A2 _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _00297_ clknet_leaf_65_clock mem.mem_dff.data_mem\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__B1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05589__I _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _00228_ clknet_leaf_102_clock mem.mem_dff.code_mem\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09234__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06048__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10567_ _00159_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10689__CLK clknet_leaf_67_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_144_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ _00090_ clknet_leaf_117_clock mem.mem_dff.code_mem\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08745__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05559__B2 _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11119_ _00711_ clknet_leaf_151_clock stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09524__I _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 i_la_addr[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10304__A1 _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10304__B2 _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06660_ _02161_ _02155_ _02151_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05611_ stack\[30\]\[7\] _01140_ _01141_ stack\[31\]\[7\] _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06591_ _02037_ _02103_ _02092_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07979__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_69_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08330_ mem.mem_dff.code_mem\[25\]\[6\] _02789_ _02846_ mem.mem_dff.code_mem\[27\]\[6\]
+ _03519_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05542_ _01042_ stack\[0\]\[6\] stack\[1\]\[6\] _01084_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08276__A3 _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09399__C _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ mem.mem_dff.code_mem\[8\]\[4\] _03292_ _03293_ mem.mem_dff.code_mem\[22\]\[4\]
+ mem.mem_dff.code_mem\[31\]\[4\] _02957_ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05473_ _01023_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__B1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05499__I _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07212_ _02597_ _02592_ _02583_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _03386_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07143_ _02543_ _02538_ _02544_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06832__B _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07074_ _02370_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__I _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05342__S0 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06025_ _01405_ _01567_ _01568_ _01476_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08736__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ _03187_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspell_264 o_wb_data[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_214_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09715_ _04480_ _04674_ single_step _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ mem.mem_dff.code_mem\[10\]\[6\] _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09646_ cycles_per_ms\[6\] _04576_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06858_ _02023_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A2 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05809_ _01330_ stack\[14\]\[0\] _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09577_ cycles_per_ms\[14\] _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ _02143_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07889__I _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08528_ _01829_ _03671_ _03686_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05630__C net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _01588_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09216__A2 _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _00013_ clknet_leaf_122_clock mem.mem_dff.code_mem\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08975__A1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__B1 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _05075_ _05153_ _05155_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05333__S0 _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05789__A1 _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ _03909_ _03232_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09775__I0 exec.memory_input\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05805__C _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05713__A1 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_70_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06269__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10619_ _00211_ clknet_leaf_105_clock mem.mem_dff.code_mem\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09758__A3 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08966__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08423__I _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06441__A2 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07039__I mem.mem_dff.code_mem\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08718__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07830_ _03079_ _03074_ _03066_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06878__I _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05782__I stack\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07941__A2 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08298__C _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _03025_ _03020_ _03026_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05952__A1 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10704__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__B2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _04441_ _04325_ _04464_ _04402_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06712_ _02102_ _02203_ _02195_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07692_ _02958_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ _04395_ _04389_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06643_ mem.mem_dff.code_mem\[3\]\[3\] _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05704__A1 _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09362_ net92 _04291_ _04292_ net83 _04306_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06574_ mem.mem_dff.code_mem\[1\]\[7\] _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10854__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08249__A3 _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08313_ _03496_ _03497_ _03502_ _03503_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05525_ _01074_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09293_ _04266_ _04276_ _04277_ _04264_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10056__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ mem.mem_dff.code_mem\[2\]\[3\] _02098_ _02588_ mem.mem_dff.code_mem\[18\]\[3\]
+ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05456_ _00921_ _01005_ _01006_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05563__S0 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ mem.mem_dff.code_mem\[15\]\[1\] _03368_ _03369_ mem.mem_dff.code_mem\[29\]\[1\]
+ mem.mem_dff.code_mem\[30\]\[1\] _02927_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05387_ stack\[6\]\[3\] _00934_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10213__B1 _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ mem.mem_dff.code_mem\[16\]\[0\] _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07057_ _02389_ _02473_ _02464_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06432__A2 _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput140 net140 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput151 net151 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08709__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput162 net162 o_wb_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06008_ stack\[30\]\[1\] stack\[31\]\[1\] _01391_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput173 net173 o_wb_data[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput184 net184 o_wb_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput195 net195 rambus_wb_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06196__A1 _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07932__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ _03167_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output136_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09134__B2 stack\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10103__I _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10970_ _00562_ clknet_leaf_43_clock net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09629_ _04583_ _04584_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06737__B _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07999__A2 _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06671__A2 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10404_ _01125_ _05188_ _05191_ stack\[15\]\[6\] _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10335_ _01857_ _05137_ _05135_ stack\[16\]\[3\] _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10266_ _05075_ _05089_ _05092_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10727__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09373__A1 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _05041_ _05042_ _05034_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10013__I _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09125__B2 stack\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09802__I _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08100__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05310_ _00789_ _00863_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06290_ _01717_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 i_wb_addr[11] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_05241_ _00789_ _00795_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput31 i_wb_addr[21] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput42 i_wb_cyc net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 i_wb_data[19] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08939__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__B2 stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput64 i_wb_data[7] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput75 io_in[6] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09061__B1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 rambus_wb_dat_i[17] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_171_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput97 rambus_wb_dat_i[27] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06414__A2 _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09980_ _01633_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ _01792_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08167__A2 _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _03819_ _03943_ _03951_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07813_ _03065_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07914__A2 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08793_ _03893_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09116__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07744_ _03009_ _03002_ _03012_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06557__B _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09414_ net257 net139 _04378_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_41_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06626_ _00759_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09419__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06350__A1 stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__I _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06350__B2 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11032__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _04324_ _04325_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06557_ _02041_ _02074_ _02066_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05888__S _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input97_I rambus_wb_dat_i[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05508_ _01036_ stack\[3\]\[5\] _01045_ stack\[2\]\[5\] _00972_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06102__A1 _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ _04260_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06488_ _02019_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08227_ mem.mem_dff.code_mem\[15\]\[3\] _03368_ _03369_ mem.mem_dff.code_mem\[29\]\[3\]
+ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05439_ _00931_ stack\[3\]\[4\] _00924_ stack\[2\]\[4\] _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08158_ _02649_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09052__B1 _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07109_ _02500_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08089_ net76 _03273_ _03274_ net127 _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08998__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A3 _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05613__B1 stack\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10120_ _01027_ _04928_ _04983_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10051_ _04917_ _04918_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05916__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05916__B2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07851__B _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07669__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10953_ _00545_ clknet_leaf_149_clock stack\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10884_ _00476_ clknet_leaf_186_clock stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__A1 _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06341__B2 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10318_ stack\[27\]\[7\] _05118_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08701__I _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10249_ _05077_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06221__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08349__S _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05790_ stack\[18\]\[0\] stack\[19\]\[0\] stack\[16\]\[0\] stack\[17\]\[0\] _01330_
+ _00844_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06580__A1 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05383__A2 stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07460_ _02790_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07052__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ exec.memory_input\[6\] _01846_ _01746_ _01169_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07391_ _02737_ _02734_ _02727_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05930__I1 stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09130_ _04054_ _04144_ _04152_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__A1 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06342_ exec.memory_input\[4\] _01846_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08085__B2 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09821__A2 _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _03755_ _04092_ _04093_ _04100_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06273_ _00981_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08012_ _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_194_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05224_ _00778_ _00771_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09034__B1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07936__B _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_192_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06938__A3 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09963_ delay_cycles\[17\] _04854_ _04852_ _04520_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08914_ _03887_ _03984_ _03969_ _03987_ _03988_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_213_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _04802_ _04701_ _04690_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07899__A1 _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _01990_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _03882_ _03871_ _03883_ _03884_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05988_ stack\[6\]\[5\] stack\[7\]\[5\] _01463_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input12_I i_la_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07727_ mem.mem_dff.data_mem\[0\]\[3\] _02992_ _02999_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10104__C1 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08312__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10422__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07658_ _02941_ _02942_ _02945_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06609_ mem.mem_dff.code_mem\[2\]\[5\] _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07589_ mem.mem_dff.code_mem\[28\]\[5\] _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05921__I1 stack\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07897__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09328_ mem.io_data_out\[3\] _04274_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08076__A1 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05509__S0 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09812__A2 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10572__CLK clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07823__A1 _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _03909_ _04109_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09025__B1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05210__I _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__B _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11152_ _00744_ clknet_leaf_176_clock stack\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05988__I1 stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10103_ _04934_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11083_ _00675_ clknet_leaf_40_clock net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10034_ _04903_ _04904_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09780__C _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08551__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ _00528_ clknet_leaf_143_clock stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06314__A1 _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10867_ _00459_ clknet_leaf_190_clock stack\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05912__I1 stack\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A1 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08067__B2 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10798_ _00390_ clknet_leaf_163_clock stack\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__A1 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06216__I _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09567__A1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10177__A2 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A1 _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06960_ _02366_ _02399_ _02395_ _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05991__S _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I i_la_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ stack\[26\]\[3\] stack\[27\]\[3\] _01410_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06891_ _02341_ _02334_ _02343_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08542__A2 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ _03696_ _03763_ _03760_ stack\[3\]\[7\] _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10445__CLK clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05842_ _01266_ _01384_ _01385_ _01290_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ _03712_ _03700_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05773_ _01015_ _01315_ _01316_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07512_ _02816_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_139_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08492_ _03656_ _03641_ _03657_ stack\[19\]\[4\] _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06305__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10595__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07443_ mem.mem_dff.code_mem\[24\]\[5\] _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06835__B _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07374_ _02641_ _02718_ _02713_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09255__B1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ net42 net67 _01626_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06325_ _01724_ net61 _01863_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09044_ _03629_ _03770_ _01616_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_136_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06256_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09558__A1 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05207_ mem.select _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09558__B2 _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06187_ _01221_ _01729_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10168__A2 _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_150_clock clknet_4_5_0_clock clknet_leaf_150_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A2 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _04819_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _04766_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08533__A2 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06796__I _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08828_ stack\[7\]\[2\] _03916_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10340__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05978__S0 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output216_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08759_ _03861_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10938__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10721_ _00313_ clknet_leaf_29_clock mem.mem_dff.data_mem\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06847__A2 _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08049__A1 _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ _00244_ clknet_leaf_94_clock mem.mem_dff.code_mem\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_103_clock clknet_4_13_0_clock clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09246__B1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ _00175_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05283__A1 _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_118_clock clknet_4_12_0_clock clknet_leaf_118_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10159__A2 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11135_ _00727_ clknet_leaf_151_clock stack\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08772__A2 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10468__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06783__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11066_ _00658_ clknet_leaf_131_clock net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10017_ delay_counter\[2\] _04648_ _04885_ _00919_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08524__A2 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09721__B2 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05824__B _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06535__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10331__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_140_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10095__A1 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10095__B2 _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _00511_ clknet_leaf_147_clock stack\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout247_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__I0 stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05510__A2 _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10398__A2 _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06110_ _01653_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07090_ _02500_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06041_ _01582_ _01584_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07486__B _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08212__A1 mem.mem_dff.code_mem\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_65_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09800_ _04729_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08763__A2 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_82_clock clknet_4_15_0_clock clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09960__B2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07992_ _03185_ _03193_ _03203_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_214_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05821__I0 stack\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06943_ _02351_ _02386_ _02378_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09731_ _03594_ _04683_ _04689_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09662_ _04621_ _04523_ _04513_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06874_ _02314_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07505__I mem.mem_dff.code_mem\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10322__A2 _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97_clock clknet_4_13_0_clock clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08613_ _03754_ _03756_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05825_ _00820_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09593_ _04550_ _04552_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08544_ _03645_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05756_ stack\[22\]\[2\] stack\[23\]\[2\] _01261_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10086__A1 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_clock clknet_4_8_0_clock clknet_leaf_20_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08475_ _03644_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05687_ _01204_ _01210_ _01226_ _01230_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_211_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05888__I0 stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07426_ _02704_ _02765_ _02756_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07240__I _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09779__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _02710_ _02705_ _02697_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_clock clknet_4_10_0_clock clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ _01026_ _01745_ _01779_ _00918_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ _02597_ _02653_ _02645_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09027_ _04004_ _04070_ _04074_ stack\[9\]\[1\] _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ exec.memory_input\[1\] _01744_ _01780_ _00841_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10610__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08203__A1 mem.mem_dff.code_mem\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output166_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09951__A1 delay_cycles\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08754__A2 _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__A2 stack\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09929_ _04556_ _04824_ _04820_ _04830_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10760__CLK clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09703__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09703__B2 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07415__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10313__A2 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11116__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10077__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _00296_ clknet_leaf_29_clock mem.mem_dff.data_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09219__B1 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08690__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10635_ _00227_ clknet_leaf_100_clock mem.mem_dff.code_mem\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _00158_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08442__A1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10497_ _00089_ clknet_leaf_117_clock mem.mem_dff.code_mem\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09077__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05559__A2 stack\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11118_ _00710_ clknet_leaf_141_clock stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11049_ _00641_ clknet_leaf_25_clock delay_cycles\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 i_la_addr[6] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10304__A2 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07325__I _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__A2 _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05610_ _01144_ stack\[28\]\[7\] stack\[29\]\[7\] _01150_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06590_ mem.mem_dff.code_mem\[2\]\[1\] _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10068__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05541_ _01086_ _01088_ _01089_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08276__A4 _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ mem.mem_dff.code_mem\[23\]\[4\] _02731_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05472_ _01000_ _01022_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08681__A1 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07060__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08681__B2 stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07211_ _02357_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ mem.dff_data_out\[1\] _03385_ _03336_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07995__I _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _02478_ _02539_ _02528_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10633__CLK clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10240__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07073_ mem.mem_dff.code_mem\[14\]\[5\] _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05729__B _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05342__S1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06024_ stack\[12\]\[1\] stack\[13\]\[1\] _01427_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10783__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07944__B _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06747__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _01683_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06926_ _02369_ _02364_ _02372_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09714_ _04648_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xspell_265 o_wb_data[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06857_ mem.mem_dff.code_mem\[9\]\[0\] _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09645_ _04588_ _04604_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ stack\[15\]\[0\] _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09576_ _04530_ _04535_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06788_ mem.mem_dff.code_mem\[7\]\[1\] _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _03654_ _03677_ _03682_ stack\[29\]\[3\] _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05739_ stack\[10\]\[2\] stack\[11\]\[2\] _00940_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08121__B1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _01604_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08672__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ mem.mem_dff.code_mem\[23\]\[6\] _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ net120 _03573_ _03576_ _03073_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10420_ _00012_ clknet_leaf_122_clock mem.mem_dff.code_mem\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__A1 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10231__A1 _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08975__A2 _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10231__B2 stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _03643_ _03996_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06986__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05333__S1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05789__A2 _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _05064_ _05097_ _05104_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__I1 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08360__B1 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09360__I _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_13_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__B1 _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10656__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08663__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05316__I2 stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08415__A1 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10618_ _00210_ clknet_leaf_105_clock mem.mem_dff.code_mem\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08704__I _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08415__B2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08966__A2 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ _00141_ clknet_leaf_76_clock mem.mem_dff.code_mem\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06977__A1 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__A2 _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ _02936_ _03021_ _03011_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06711_ _02201_ _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10289__A1 _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07691_ mem.mem_dff.code_mem\[31\]\[4\] _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08351__B1 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09430_ _04402_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06642_ _02146_ _02139_ _02147_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06901__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09361_ net106 _04304_ _02134_ net101 _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06573_ _02089_ _02084_ _02090_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ mem.mem_dff.code_mem\[11\]\[5\] _03299_ _02414_ mem.mem_dff.code_mem\[12\]\[5\]
+ mem.mem_dff.code_mem\[26\]\[5\] _03300_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05524_ _01073_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _03622_ _01727_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10056__A4 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05303__I _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08243_ mem.mem_dff.code_mem\[5\]\[3\] _02200_ _02650_ mem.mem_dff.code_mem\[20\]\[3\]
+ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05455_ _00931_ stack\[19\]\[4\] _00933_ stack\[18\]\[4\] _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05563__S1 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07209__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _02901_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08406__A1 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__B2 _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05386_ _00937_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07125_ _02525_ _02516_ _02529_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10213__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10213__B2 stack\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08421__A4 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07056_ mem.mem_dff.code_mem\[14\]\[1\] _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06134__I _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput130 net130 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput141 net141 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09906__A1 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 net152 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06007_ _01409_ _01549_ _01550_ _01414_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput163 net163 o_wb_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput174 net174 o_wb_data[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput185 net185 rambus_wb_addr_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input42_I i_wb_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09445__I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput196 net196 rambus_wb_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10529__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06196__A2 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07958_ _02996_ _03171_ _03175_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05943__A2 stack\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09134__A2 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06909_ _02358_ _02352_ _02342_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output129_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ _01998_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08342__B1 _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10679__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09628_ cycles_per_ms\[4\] _04582_ _04586_ _04587_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ cycles_per_ms\[17\] _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_187_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05213__I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10403_ _05183_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09070__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10334_ _05057_ _05141_ _05143_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06044__I _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05482__I1 stack\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06979__I _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _05092_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08176__A3 _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09373__A2 mem.dff_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ _04500_ _05032_ _05037_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07384__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05395__B1 _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09125__A2 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07136__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08884__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05698__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05551__C _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06219__I _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05240_ stack\[3\]\[0\] stack\[0\]\[0\] stack\[1\]\[0\] stack\[2\]\[0\] _00792_ _00794_
+ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08434__I _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 i_la_data[2] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_204_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput21 i_wb_addr[12] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput32 i_wb_addr[22] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 i_wb_data[0] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08939__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 i_wb_data[1] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09061__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput65 i_wb_data[8] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput76 io_in[7] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09061__B2 _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05994__S _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput87 rambus_wb_dat_i[18] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput98 rambus_wb_dat_i[28] net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ _03992_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06889__I _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08861_ _03776_ _03947_ _03950_ stack\[26\]\[0\] _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07812_ _01998_ _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08792_ _03207_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10821__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09116__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ mem.mem_dff.data_mem\[0\]\[7\] _03003_ _03011_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__B1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07674_ _02874_ _02957_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08875__A1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06625_ net255 _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09413_ _04387_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10971__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06350__A2 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06556_ mem.mem_dff.code_mem\[1\]\[2\] _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08627__A1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09344_ _01864_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05507_ _01049_ _01056_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_205_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09275_ _01662_ _01663_ _01664_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_205_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07669__B _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06487_ net255 _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08226_ _03419_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05438_ _00923_ _00988_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08157_ _02199_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09052__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05369_ _00887_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09052__B2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _02500_ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _03282_ _03285_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10201__A4 _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05613__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07039_ mem.mem_dff.code_mem\[13\]\[6\] _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05613__B2 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09355__A2 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10050_ net41 net40 net20 net19 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_130_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05377__B1 stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09903__I _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07118__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10952_ _00544_ clknet_leaf_144_clock stack\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _00475_ clknet_leaf_193_clock stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06341__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06039__I _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09778__C _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05878__I _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05852__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05604__A1 stack\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _05066_ _05129_ _05130_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05604__B2 stack\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10844__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09346__A2 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _05057_ _05072_ _05081_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05546__C _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07357__A1 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ net170 _05023_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10361__B1 _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09813__I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06580__A2 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _01801_ _01945_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07390_ _02505_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05391__I0 stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06341_ _01859_ _01808_ _01877_ _01878_ _01879_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__A2 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _00919_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08164__I _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ _01795_ _01808_ _01810_ _01579_ _01812_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_191_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ _01855_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05223_ net140 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09034__B2 stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08242__C1 mem.mem_dff.code_mem\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_135_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06938__A4 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _04823_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08913_ stack\[10\]\[7\] _03976_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06412__I _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09893_ _04678_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _03846_ _03934_ _03935_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08775_ stack\[11\]\[5\] _03862_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05987_ stack\[4\]\[5\] stack\[5\]\[5\] _01442_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07726_ _02952_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ _02943_ _02944_ _02939_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07520__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05899__S _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06608_ _02114_ _02115_ _02119_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ _02888_ _02889_ _02891_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10407__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10717__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06539_ _02063_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09327_ _04268_ mem.dff_data_out\[3\] _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05509__S1 _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__A1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08074__I _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _04180_ _04233_ _04245_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05834__A1 _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08209_ mem.mem_dff.code_mem\[5\]\[2\] _02200_ _02650_ mem.mem_dff.code_mem\[20\]\[2\]
+ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09189_ _04122_ _04192_ _04189_ stack\[20\]\[1\] _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09025__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09025__B2 stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10867__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11151_ _00743_ clknet_4_7_0_clock stack\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05598__B1 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10102_ net177 _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11082_ _00674_ clknet_leaf_125_clock delay_counter\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06322__I _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10033_ delay_counter\[5\] _04674_ _04899_ _01075_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_1_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10343__B1 _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08551__A3 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08839__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07153__I mem.mem_dff.code_mem\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09500__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ _00527_ clknet_leaf_143_clock stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ _00458_ clknet_leaf_183_clock stack\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10797_ _00389_ clknet_leaf_134_clock stack\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05401__I _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07578__A1 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08378__I0 mem.dff_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ _01355_ _01450_ _01453_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06890_ _02282_ _02335_ _02342_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ stack\[14\]\[7\] stack\[15\]\[7\] _01013_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05772_ _01264_ stack\[30\]\[2\] _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08560_ _01795_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07511_ _02050_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08491_ _03647_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__I _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_61_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ _02774_ _02775_ _02777_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ mem.mem_dff.code_mem\[22\]\[6\] _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__B2 stack\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06069__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _04137_ _04134_ _04114_ _04112_ _04138_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06324_ _01721_ _01862_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09270__A4 _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09043_ _03636_ _01685_ _01930_ _03663_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06255_ _01795_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05206_ _00762_ net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06186_ _01728_ _01210_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13_0_clock clknet_3_6_0_clock clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07569__A1 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10092__C _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__A1 _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06142__I _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _04840_ _04842_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09876_ _03281_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__B1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08827_ _03922_ _03923_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__B _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05978__S1 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _03870_ _03824_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output111_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07709_ net254 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output209_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03791_ _03809_ _03814_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10720_ _00312_ clknet_leaf_31_clock mem.mem_dff.data_mem\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _00243_ clknet_leaf_94_clock mem.mem_dff.code_mem\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09246__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09246__B2 stack\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10582_ _00174_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06317__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11045__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11134_ _00726_ clknet_leaf_145_clock stack\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11065_ _00657_ clknet_leaf_20_clock delay_cycles\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_49_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10316__B1 _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05418__S0 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _04880_ _04886_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09721__A2 _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08288__A2 _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09485__A1 _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06299__A1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10918_ _00510_ clknet_leaf_148_clock stack\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07611__I mem.mem_dff.code_mem\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09237__A1 stack\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05897__I1 stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10849_ _00441_ clknet_leaf_162_clock stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__B1 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06040_ _01321_ _01240_ _01583_ _00778_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_201_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10412__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09960__A2 _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _03198_ _03202_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09730_ _04658_ _04684_ _04688_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__05821__I1 stack\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06942_ _02384_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10307__B1 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09661_ _04507_ _04508_ _04520_ _04519_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06873_ mem.mem_dff.code_mem\[9\]\[3\] _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08612_ _03755_ _03748_ _03749_ net146 _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_209_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05824_ _01291_ _01364_ _01278_ _01367_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09592_ _04551_ _04547_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05755_ _01298_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08543_ _01991_ _03693_ _03697_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08279__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10086__A2 _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input107_I rambus_wb_dat_i[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08474_ _03628_ _03199_ _01636_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05686_ _01189_ _01229_ _01213_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07425_ _02763_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05888__I1 stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09779__A2 _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07356_ _02357_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11068__CLK clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06307_ exec.memory_input\[3\] _01846_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ mem.mem_dff.code_mem\[20\]\[2\] _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07677__B _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input72_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09026_ _04066_ _04068_ _04075_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06238_ _01779_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06169_ _01704_ _01711_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_172_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output159_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06765__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__CLK clknet_leaf_181_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _04573_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09183__I _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A2 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _04610_ _04769_ _04780_ net45 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09911__I _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10703_ _00295_ clknet_leaf_66_clock mem.mem_dff.data_mem\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09219__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09219__B2 stack\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08690__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10634_ _00226_ clknet_leaf_101_clock mem.mem_dff.code_mem\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10565_ _00157_ clknet_leaf_73_clock mem.mem_dff.code_mem\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05886__I _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06453__A1 _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06453__B2 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10496_ _00088_ clknet_leaf_116_clock mem.mem_dff.code_mem\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10001__A2 _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A3 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07953__A1 mem.mem_dff.data_mem\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11117_ _00709_ clknet_leaf_141_clock stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11048_ _00640_ clknet_leaf_26_clock delay_cycles\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 i_la_data[0] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08902__B1 _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06666__B _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05540_ _00920_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05471_ _00854_ _01008_ _01021_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08681__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07210_ mem.mem_dff.code_mem\[18\]\[2\] _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06692__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08190_ _03374_ _03384_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07141_ mem.mem_dff.code_mem\[16\]\[2\] _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08969__B1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06444__A1 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07072_ _02483_ _02484_ _02487_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10240__A2 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10928__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06023_ stack\[14\]\[1\] stack\[15\]\[1\] _00810_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_179_clock clknet_4_4_0_clock clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ _01675_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_clock clknet_4_13_0_clock clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09713_ _04286_ _04667_ _04669_ _04672_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06925_ _02371_ _02367_ _02361_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xspell_266 o_wb_data[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09697__A1 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07960__B _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ _04603_ _04590_ _04581_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06856_ _02313_ _02306_ _02316_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05807_ stack\[12\]\[0\] stack\[13\]\[0\] _01330_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09575_ delay_cycles\[13\] _04534_ delay_cycles\[14\] _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06787_ _02254_ _02260_ _02262_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_clock clknet_4_12_0_clock clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08526_ _01797_ _03671_ _03685_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05738_ _01281_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08457_ _03619_ _03624_ _03626_ _03627_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08672__A2 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05669_ _01211_ _01212_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__CLK clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__A1 _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07408_ _02749_ _02746_ _02750_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08388_ _03575_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ mem.mem_dff.code_mem\[21\]\[7\] _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A1 _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10231__A2 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _05153_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06986__A2 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _04013_ _04043_ _04057_ stack\[25\]\[5\] _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10281_ _01923_ _05089_ _05101_ stack\[30\]\[5\] _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_183_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05797__I0 stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_207_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__A1 mem.mem_dff.code_mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07161__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_clock clknet_4_15_0_clock clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09860__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05316__I3 stack\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06674__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _00209_ clknet_leaf_106_clock mem.mem_dff.code_mem\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06505__I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _00140_ clknet_leaf_76_clock mem.mem_dff.code_mem\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_96_clock clknet_4_15_0_clock clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05549__C _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06977__A2 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10479_ _00071_ clknet_leaf_114_clock mem.mem_dff.code_mem\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__I _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07926__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07336__I mem.mem_dff.code_mem\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06240__I _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09679__A1 _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06710_ _02201_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07690_ _02967_ _02959_ _02970_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_34_clock clknet_4_8_0_clock clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08351__A1 mem.mem_dff.code_mem\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08351__B2 mem.mem_dff.code_mem\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06641_ _02109_ _02140_ _02130_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09360_ _04338_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06572_ _02060_ _02085_ _02081_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10600__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08311_ _03498_ _03499_ _03500_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05523_ _01072_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49_clock clknet_4_11_0_clock clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09291_ _04267_ _04273_ _04275_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08242_ mem.mem_dff.code_mem\[3\]\[3\] _02137_ _02173_ mem.mem_dff.code_mem\[4\]\[3\]
+ mem.mem_dff.code_mem\[21\]\[3\] _02676_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05454_ _00924_ _01004_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10750__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ _02498_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05385_ _00799_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07124_ _02527_ _02517_ _02528_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10213__A2 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07055_ _02466_ _02471_ _02474_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07955__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput120 net120 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput131 net131 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__11106__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06006_ stack\[24\]\[1\] stack\[25\]\[1\] _01329_ _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput142 net256 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput153 net153 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput164 net164 o_wb_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput175 net175 o_wb_data[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07917__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput186 net254 rambus_wb_addr_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput197 net197 rambus_wb_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05779__I0 stack\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__I mem.mem_dff.code_mem\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input35_I i_wb_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07957_ mem.mem_dff.data_mem\[7\]\[2\] _03172_ _03168_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07888_ _02063_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08342__B2 _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ cycles_per_ms\[3\] _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06839_ _02269_ _02296_ _02303_ _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08893__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09558_ _04514_ _04495_ _04515_ _04516_ _04517_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_102_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05951__I0 stack\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08509_ _03670_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09842__A1 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _01667_ _04299_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10402_ _05190_ _05192_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09070__A2 _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _01825_ _05137_ _05135_ stack\[16\]\[2\] _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07865__B _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05631__A2 _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05482__I2 stack\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _01638_ _03198_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10195_ net175 _05035_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07156__I mem.mem_dff.code_mem\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08581__A1 stack\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06060__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05395__A1 stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05395__B2 _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10623__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10140__A1 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05698__A2 _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10773__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09833__A1 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06647__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 i_la_data[3] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput22 i_wb_addr[13] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11129__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 i_wb_addr[23] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 i_wb_data[10] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput55 i_wb_data[20] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput66 i_wb_data[9] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__09061__A2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput77 rambus_wb_ack_i net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput88 rambus_wb_dat_i[19] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 rambus_wb_dat_i[29] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09349__B1 _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08450__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08860_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__B _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08572__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ mem.mem_dff.data_mem\[2\]\[7\] _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ stack\[6\]\[0\] _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_211_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ _03010_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09281__I _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08324__A1 mem.mem_dff.code_mem\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05515__S _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08875__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10131__B2 _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_131_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09412_ _04338_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06624_ mem.mem_dff.code_mem\[3\]\[0\] _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06886__A1 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06555_ _02076_ _02073_ _02077_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08627__A2 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06638__A1 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05506_ _01030_ stack\[0\]\[5\] stack\[1\]\[5\] _01031_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09274_ _03620_ _04258_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06486_ _02017_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ mem.dff_data_out\[2\] _03418_ _03336_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05437_ _00945_ stack\[0\]\[4\] stack\[1\]\[4\] _00944_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08156_ mem.mem_dff.code_mem\[2\]\[1\] _03349_ _03350_ mem.mem_dff.code_mem\[18\]\[1\]
+ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05368_ _00908_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A1 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09052__A2 _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07107_ mem.mem_dff.code_mem\[15\]\[4\] _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ mem.io_data_out\[6\] _03267_ _03271_ _03284_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05299_ _00850_ _00772_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__A1 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05613__A2 stack\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07038_ _02459_ _02456_ _02460_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_56_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05917__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10646__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08563__A1 _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output141_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05377__A1 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ stack\[25\]\[0\] _04046_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05377__B2 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10370__A1 stack\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07704__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08315__B2 mem.mem_dff.data_mem\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _00543_ clknet_leaf_143_clock stack\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10796__CLK clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10122__A1 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10882_ _00474_ clknet_leaf_183_clock stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__B1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09815__A1 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_3_0_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07054__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10316_ _05068_ _05115_ _05118_ stack\[27\]\[6\] _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _04220_ _05074_ _05078_ stack\[14\]\[2\] _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08554__A1 _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10178_ _05027_ _05028_ _05022_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10361__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08306__A1 mem.mem_dff.code_mem\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08306__B2 mem.mem_dff.code_mem\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07614__I mem.mem_dff.code_mem\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05335__S _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10113__A1 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05562__C _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06868__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08609__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06340_ _01023_ _01878_ _01809_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_206_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08445__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10519__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06271_ _00918_ _01811_ _01579_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_198_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05222_ net140 _00776_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08010_ _01797_ _03213_ _03219_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05843__A2 _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09034__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__C2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10669__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09961_ _04850_ _04853_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05446__I2 stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _03855_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10215__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09892_ _04799_ _04801_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09742__B1 _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03851_ _03930_ _03928_ stack\[7\]\[6\] _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__A1 _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ _03228_ _03859_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05986_ _01259_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07524__I _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ _02149_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__A1 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__B2 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07656_ _02928_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06607_ _02117_ _02118_ _02112_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07587_ _02831_ _02890_ _02886_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ _04305_ _04307_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06538_ net233 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06087__A2 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__B _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _04227_ _04235_ _04242_ stack\[22\]\[5\] _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06469_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ mem.mem_dff.code_mem\[3\]\[2\] _02137_ _02173_ mem.mem_dff.code_mem\[4\]\[2\]
+ mem.mem_dff.code_mem\[21\]\[2\] _02676_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_182_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09025__A2 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output189_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ _02014_ _03334_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06603__I _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11150_ _00742_ clknet_leaf_138_clock stack\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05598__A1 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05598__B2 stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10101_ _04966_ _04967_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11081_ _00673_ clknet_leaf_127_clock delay_counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05219__I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09914__I _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10032_ _04894_ _04895_ _04900_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10343__A1 _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10343__B2 stack\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06011__A2 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05770__A1 _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08839__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10934_ _00526_ clknet_leaf_143_clock stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10865_ _00457_ clknet_leaf_150_clock stack\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05522__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10796_ _00388_ clknet_4_0_0_clock stack\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10811__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10961__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08378__I1 _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__B2 stack\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10334__A1 _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05840_ stack\[12\]\[7\] stack\[13\]\[7\] _00770_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05771_ stack\[31\]\[2\] _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05761__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07510_ _02816_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08490_ _03223_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _02717_ _02776_ _02772_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05513__A1 stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07372_ _02720_ _02716_ _02722_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09255__A2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ stack\[24\]\[7\] _04120_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06323_ net12 _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06069__A2 _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10491__CLK clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _04019_ _04082_ _04067_ _03987_ _04084_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06254_ _00916_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05205_ _00756_ mem.addr\[0\] _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08215__B1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09558__A3 _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06185_ _01578_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07569__A2 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07519__I mem.mem_dff.code_mem\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05467__C _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09944_ _04544_ _04835_ _04832_ _04841_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08518__A1 _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09875_ _04784_ _04790_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__B2 stack\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ _03215_ _03919_ _03920_ net145 _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07254__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08757_ _03645_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05969_ _01505_ _01512_ _01446_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ _02101_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08688_ _03656_ _03800_ _03813_ stack\[5\]\[4\] _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09494__A2 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ _02928_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05504__A1 _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10650_ _00242_ clknet_leaf_101_clock mem.mem_dff.code_mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10834__CLK clknet_leaf_177_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09246__A2 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09309_ _00762_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _00173_ clknet_leaf_84_clock mem.mem_dff.code_mem\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07009__A1 _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08206__B1 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10984__CLK clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09954__B1 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11133_ _00725_ clknet_leaf_152_clock stack\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06232__A2 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07873__B _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05291__I0 stack\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11064_ _00656_ clknet_leaf_21_clock delay_cycles\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10316__A1 _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10316__B2 stack\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10015_ _04884_ _04887_ _04889_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05418__S1 _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07164__I mem.mem_dff.code_mem\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05743__A1 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05743__B2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07496__A1 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ _00509_ clknet_leaf_147_clock stack\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_178_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__B1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10848_ _00440_ clknet_leaf_161_clock stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09237__A2 _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07248__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10779_ _00371_ clknet_leaf_41_clock mem.io_data_ready vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10252__B1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__B2 stack\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07990_ _03201_ _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06941_ _02384_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10307__A1 _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10707__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__B2 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__A1 _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05982__B2 _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__A1 _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ _04571_ _04609_ _04615_ _04616_ _04617_ _04619_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_67_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06872_ _02328_ _02323_ _02329_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07074__I _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ _03217_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05823_ _01303_ _01365_ _01366_ _01290_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09591_ cycles_per_ms\[12\] _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _03696_ _03680_ _03687_ stack\[29\]\[7\] _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05754_ _01280_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10857__CLK clknet_leaf_168_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09476__A2 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08473_ _03629_ _03194_ _03195_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05685_ _01227_ _01228_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__B1 stack\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07424_ _02763_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05322__I _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07355_ mem.mem_dff.code_mem\[22\]\[2\] _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__B1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06306_ _01246_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08633__I _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ _02655_ _02652_ _02656_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09025_ _04024_ _04070_ _04074_ stack\[9\]\[0\] _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06237_ _01248_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input65_I i_wb_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07411__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06099_ net110 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ _04798_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05973__A1 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05973__B2 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10403__I _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _04774_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07714__A2 _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08911__A1 _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output221_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08809_ _01713_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09789_ _04723_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05725__A1 _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08808__I _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _00294_ clknet_leaf_66_clock mem.mem_dff.data_mem\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09219__A2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11012__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _00225_ clknet_leaf_101_clock mem.mem_dff.code_mem\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07868__B _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10564_ _00156_ clknet_leaf_82_clock mem.mem_dff.code_mem\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10495_ _00087_ clknet_leaf_117_clock mem.mem_dff.code_mem\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07159__I mem.mem_dff.code_mem\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11162__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__A4 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11116_ _00708_ clknet_leaf_141_clock stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05964__A1 _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05964__B2 _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11047_ _00639_ clknet_leaf_26_clock delay_cycles\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06012__B _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08902__A1 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 i_la_data[1] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08902__B2 stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06947__B _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05570__C _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__B1 _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10068__A3 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08130__A2 _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05470_ _01017_ _01018_ _01020_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08969__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ _02541_ _02538_ _02542_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08969__B2 stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07071_ _02485_ _02486_ _02481_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07069__I _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09769__I0 exec.memory_input\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06022_ _01011_ _01564_ _01565_ _01286_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06701__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07973_ _02002_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05955__A1 _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09146__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ _04670_ _04671_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06924_ _02370_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspell_267 rambus_wb_addr_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09697__A2 _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ cycles_per_ms\[2\] _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06855_ _02282_ _02307_ _02315_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05806_ _00944_ _01346_ _01349_ _01313_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09574_ _04532_ delay_cycles\[11\] delay_cycles\[10\] _04533_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06786_ _02229_ _02261_ _02252_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06380__B2 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _03652_ _03677_ _03682_ stack\[29\]\[2\] _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05737_ _01280_ _01265_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _03568_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06148__I _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06132__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05668_ net158 _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08672__A3 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07407_ _02721_ _02747_ _02743_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08387_ mem.mem_io.past_write _03574_ _03570_ _03571_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_05599_ _01129_ _01145_ _01146_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10216__B1 _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07338_ _02694_ _02689_ _02695_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09621__A2 _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06435__A2 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _02640_ _02635_ _02642_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _01892_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output171_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10280_ _05061_ _05098_ _05103_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__A2 _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_clock clknet_4_0_0_clock clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06611__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05946__A1 _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05797__I1 stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09137__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10133__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05961__A4 _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08360__A2 _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__I _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06371__A1 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__A2 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06123__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07598__B _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10616_ _00208_ clknet_leaf_105_clock mem.mem_dff.code_mem\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05309__S0 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10552__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _00139_ clknet_leaf_79_clock mem.mem_dff.code_mem\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06977__A3 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10478_ _00070_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06521__I _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05937__A1 _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10289__A3 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06677__B _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08351__A2 _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06640_ mem.mem_dff.code_mem\[3\]\[2\] _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06362__A1 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07352__I mem.mem_dff.code_mem\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06571_ mem.mem_dff.code_mem\[1\]\[6\] _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08310_ mem.mem_dff.code_mem\[3\]\[5\] _03364_ _03365_ mem.mem_dff.code_mem\[4\]\[5\]
+ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09300__A1 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05522_ _00979_ _01055_ _01071_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ mem.io_data_out\[0\] _04274_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06114__A1 _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _03424_ _03427_ _03431_ _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05453_ _00945_ stack\[16\]\[4\] stack\[17\]\[4\] _00962_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09500__C _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09279__I _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ mem.mem_dff.code_mem\[3\]\[1\] _03364_ _03365_ mem.mem_dff.code_mem\[4\]\[1\]
+ mem.mem_dff.code_mem\[19\]\[1\] _03366_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08183__I _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05384_ _00922_ _00930_ _00935_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07123_ _02494_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10218__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07054_ _02472_ _02473_ _02464_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput121 net121 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput132 net132 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_217_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09367__A1 _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06005_ stack\[26\]\[1\] stack\[27\]\[1\] _01412_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput143 net143 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput154 net154 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput165 net165 o_wb_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput176 net176 o_wb_data[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07917__A2 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 net187 rambus_wb_addr_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput198 net198 rambus_wb_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07971__B _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ _02994_ _03171_ _03174_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I i_wb_addr[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ net244 _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ mem.mem_dff.data_mem\[4\]\[7\] _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06838_ _02251_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09626_ delay_cycles\[3\] _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08893__A3 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09557_ cycles_per_ms\[18\] _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06769_ _02245_ _02241_ _02247_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05951__I1 stack\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08508_ _03198_ _03669_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_197_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09488_ _01130_ _04449_ _04455_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_200_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09842__A2 _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10575__CLK clknet_leaf_89_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08439_ _02056_ _03609_ _03613_ _03612_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09410__C _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06606__I _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ net149 _05188_ _05191_ stack\[15\]\[5\] _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10128__I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08802__B1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10332_ _05053_ _05141_ _05142_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08821__I _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05631__A3 _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10263_ _03898_ _05090_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08030__A1 _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _05039_ _05040_ _05034_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08581__A2 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07881__B _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05395__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_163_clock clknet_4_6_0_clock clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08333__A2 _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05698__A3 _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10918__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_178_clock clknet_4_4_0_clock clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09320__C _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__I _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06516__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_101_clock clknet_4_13_0_clock clknet_leaf_101_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 i_la_data[4] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05420__I _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 i_wb_addr[14] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput34 i_wb_addr[2] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput45 i_wb_data[11] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput56 i_wb_data[21] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput67 i_wb_stb net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05607__B1 _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput78 rambus_wb_dat_i[0] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput89 rambus_wb_dat_i[1] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08731__I _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09349__A1 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_clock clknet_4_12_0_clock clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09349__B2 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07347__I _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06251__I _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _03062_ _03057_ _03063_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07791__B _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08572__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10448__CLK clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06583__A1 _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07741_ _02840_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07672_ _02787_ _02412_ _02255_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_26_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06335__A1 _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10131__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06335__B2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ net257 _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06623_ _02126_ _02115_ _02131_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10598__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05933__I1 stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _03620_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06554_ _02037_ _02074_ _02066_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05505_ _01039_ _01054_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09273_ _04249_ _04257_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06485_ _02016_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08224_ _03412_ _03417_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05436_ stack\[6\]\[4\] _00984_ _00959_ stack\[7\]\[4\] _00921_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06426__I _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05330__I _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08155_ _02587_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09588__B2 cycles_per_ms\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07966__B _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05367_ _00919_ net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07106_ _02510_ _02501_ _02514_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08641__I _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__A1 mem.mem_dff.code_mem\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ net118 _03272_ _03283_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05298_ _00851_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07037_ _02371_ _02457_ _02453_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_clock clknet_4_15_0_clock clknet_leaf_80_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08563__A2 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08988_ _04045_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05377__A2 stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10370__A2 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output134_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07939_ _03154_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10950_ _00542_ clknet_leaf_144_clock stack\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_clock clknet_4_15_0_clock clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _04564_ _04566_ _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10881_ _00473_ clknet_leaf_179_clock stack\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05924__I1 stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__A1 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__B2 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_33_clock clknet_4_10_0_clock clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10315_ _03663_ _03964_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05860__I0 stack\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06071__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _05053_ _05072_ _05080_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48_clock clknet_4_9_0_clock clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08554__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10177_ _04514_ _05020_ _05025_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09382__I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05999__S0 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10361__A2 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05843__C _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10740__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08306__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05915__I1 stack\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10890__CLK clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07630__I _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07817__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06270_ _01785_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05221_ _00773_ _00774_ _00775_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07045__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09990__A1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _04509_ _04846_ _04852_ _04521_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05446__I3 stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07077__I mem.mem_dff.code_mem\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08911_ _03963_ _03984_ _03985_ _03986_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09891_ _04483_ _04768_ _04795_ net58 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09742__A1 _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09742__B2 _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _03664_ _03796_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__I mem.mem_dff.data_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08773_ _03728_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05985_ stack\[2\]\[5\] stack\[3\]\[5\] stack\[0\]\[5\] stack\[1\]\[5\] _01371_ _00869_
+ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07724_ _02996_ _02991_ _02997_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06308__A1 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06308__B2 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07655_ _02050_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06865__B _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06606_ _02099_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07586_ _02877_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08636__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ net88 _04291_ _04292_ net80 _04306_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06537_ mem.mem_dff.code_mem\[0\]\[7\] _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I rambus_wb_dat_i[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09256_ _04177_ _04233_ _04244_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06468_ _01643_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08207_ _03395_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05419_ _00938_ _00970_ _00908_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ _04193_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06399_ _01121_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10613__CLK clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08138_ _01995_ _01996_ _02008_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08069_ mem.io_data_out\[3\] _03267_ _03246_ _03269_ _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05598__A2 stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10100_ net172 _04957_ _04429_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11080_ _00672_ clknet_leaf_125_clock delay_counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10763__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _04902_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09416__B _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10343__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05235__I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10933_ _00525_ clknet_leaf_0_clock stack\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ _00456_ clknet_leaf_150_clock stack\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08546__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07450__I _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _00387_ clknet_leaf_5_clock stack\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05905__S0 _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08281__I _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08224__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08775__A2 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06786__A1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10229_ _03847_ _04016_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10334__A2 _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05770_ _00954_ _01309_ _01312_ _01313_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05761__A2 _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07440_ _02763_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08456__I _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07360__I _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05513__A2 _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _02721_ _02718_ _02713_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_99_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09110_ _03853_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10636__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06322_ _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ stack\[9\]\[7\] _04074_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06253_ _01764_ _01642_ _01794_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05204_ _00761_ net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_159_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06184_ _01722_ net43 _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10786__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10022__B2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08766__A2 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04611_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09715__A1 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ _04514_ _04785_ _04788_ net51 _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08825_ stack\[7\]\[1\] _03916_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08756_ _03868_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05968_ _01282_ _01508_ _01511_ _01307_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I i_la_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _02980_ _02972_ _02983_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05899_ stack\[6\]\[6\] stack\[7\]\[6\] _01442_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08687_ _03802_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08151__B1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__I0 stack\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ _02030_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07569_ _02874_ _02876_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _00761_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10580_ _00172_ clknet_leaf_86_clock mem.mem_dff.code_mem\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_7_0_clock clknet_3_3_0_clock clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10261__A1 _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _01715_ _04086_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06614__I mem.mem_dff.code_mem\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__A1 mem.mem_dff.code_mem\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06217__B1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ net193 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06768__A1 _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _00724_ clknet_leaf_153_clock stack\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05440__A1 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11063_ _00655_ clknet_leaf_21_clock delay_cycles\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10316__A2 _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10014_ delay_counter\[1\] _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10509__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06940__A1 _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11091__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10916_ _00508_ clknet_leaf_188_clock stack\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08693__B2 stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10847_ _00439_ clknet_leaf_161_clock stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _00370_ clknet_leaf_122_clock net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__B1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10252__B2 stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08996__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06524__I _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__B2 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06940_ _02286_ _02383_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I i_la_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10307__A2 _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ _02235_ _02324_ _02315_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08610_ stack\[3\]\[2\] _03746_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ stack\[22\]\[7\] stack\[23\]\[7\] _01013_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09590_ cycles_per_ms\[14\] _04530_ _04535_ _04543_ cycles_per_ms\[13\] _04550_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05753_ _01260_ _01296_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08541_ _01170_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09503__C _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__I _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__A1 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05684_ _01192_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07090__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _02759_ _02762_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05498__A1 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05498__B2 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _02707_ _02703_ _02708_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__A2 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10243__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06305_ _01835_ _01839_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_206_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10243__B2 stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08987__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ _02626_ _02653_ _02645_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06998__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09024_ _04073_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06236_ _01770_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06167_ _01689_ _01706_ _01708_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input58_I i_wb_data[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06098_ _01641_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09926_ _04816_ _04828_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09857_ _04779_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _01963_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09788_ _04729_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10801__CLK clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03853_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_122_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06609__I mem.mem_dff.code_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__I _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _00293_ clknet_leaf_66_clock mem.mem_dff.data_mem\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10951__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06150__A2 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08427__A1 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10632_ _00224_ clknet_leaf_115_clock mem.mem_dff.code_mem\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10234__A1 _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _00155_ clknet_4_15_0_clock mem.mem_dff.code_mem\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__A1 _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ _00086_ clknet_leaf_120_clock mem.mem_dff.code_mem\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05661__A1 _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05413__A1 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11115_ _00707_ clknet_leaf_192_clock stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11046_ _00638_ clknet_leaf_26_clock delay_cycles\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08363__B1 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08902__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06913__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08115__B1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07124__B _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08666__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09863__B1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08666__B2 stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__A1 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08418__B2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08969__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07070_ _02470_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06254__I _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06021_ stack\[8\]\[1\] stack\[9\]\[1\] _01442_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09769__I1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__B _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05404__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07972_ _03009_ _03178_ _03184_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05955__A2 stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10824__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _04276_ _04297_ _04311_ _04344_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09146__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06923_ net238 _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07157__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspell_268 rambus_wb_addr_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09642_ _04597_ _04599_ _04601_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06854_ _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06904__A1 _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05805_ _01261_ _01347_ _01348_ _00844_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06785_ _02259_ _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09573_ _04491_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08106__B1 _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05736_ _01270_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08524_ _01764_ _03671_ _03684_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__B1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05667_ net159 _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08455_ _03625_ _01243_ intr\[1\] _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_212_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ mem.mem_dff.code_mem\[23\]\[5\] _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08409__A1 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08386_ _03251_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05598_ _01087_ stack\[11\]\[7\] _01105_ stack\[10\]\[7\] _01040_ _01146_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10216__A1 _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _02641_ _02690_ _02686_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10216__B2 stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05891__A1 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05891__B2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__A1 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _02641_ _02636_ _02632_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05643__A1 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09909__A1 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ _04059_ _04052_ _04060_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06219_ _00874_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07199_ _02096_ _02586_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08188__A3 _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06113__B net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09137__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09909_ _04799_ _04815_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_219_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08896__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05444__S _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10615_ _00207_ clknet_leaf_106_clock mem.mem_dff.code_mem\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05309__S1 _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06074__I _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10546_ _00138_ clknet_leaf_79_clock mem.mem_dff.code_mem\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_4_0_clock clknet_2_2_0_clock clknet_3_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_10_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05634__A1 edge_interrupts vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10477_ _00069_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09385__I _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10847__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07387__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09128__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07139__A1 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08336__B1 _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _00621_ clknet_leaf_14_clock cycles_per_ms\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08887__A1 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10289__A4 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ _02087_ _02084_ _02088_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05521_ _00979_ _01070_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07311__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06114__A2 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ mem.mem_dff.code_mem\[12\]\[3\] _02415_ _03432_ mem.mem_dff.code_mem\[14\]\[3\]
+ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05452_ stack\[22\]\[4\] _00984_ _00993_ stack\[23\]\[4\] _01002_ _01003_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08171_ _02619_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05383_ _00932_ stack\[3\]\[3\] _00934_ stack\[2\]\[3\] _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07122_ _02526_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08811__A1 stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07053_ _02470_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput111 net111 interrupt vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput122 net122 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06004_ _01275_ _01544_ _01547_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09367__A2 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput133 net133 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput144 net144 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput155 net155 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput166 net166 o_wb_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput177 net177 o_wb_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput188 net188 rambus_wb_addr_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput199 net199 rambus_wb_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07955_ mem.mem_dff.data_mem\[7\]\[1\] _03172_ _03168_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11002__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06868__B _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06906_ mem.mem_dff.code_mem\[10\]\[2\] _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08878__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__I _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__B1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _03121_ _03116_ _03123_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09625_ delay_cycles\[2\] _04583_ _04584_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06837_ mem.mem_dff.code_mem\[8\]\[3\] _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09556_ _04485_ _04494_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11152__CLK clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06768_ _02246_ _02243_ _02238_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08507_ _03668_ _01637_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05719_ _00941_ stack\[5\]\[2\] _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06699_ _02191_ _02186_ _02192_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09487_ _02000_ _04454_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08438_ net117 _03610_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08369_ mem.mem_dff.code_mem\[11\]\[7\] _02382_ _02442_ mem.mem_dff.code_mem\[13\]\[7\]
+ mem.mem_dff.code_mem\[26\]\[7\] _02814_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10400_ _04374_ _05183_ _05169_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08802__A1 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10331_ _01793_ _05137_ _05135_ stack\[16\]\[1\] _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10262_ _05089_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _04505_ _05032_ _05037_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08030__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06592__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10125__B1 _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07541__A1 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08284__I _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09046__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 i_la_data[5] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput24 i_wb_addr[15] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 i_wb_addr[3] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput46 i_wb_data[12] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput57 i_wb_data[22] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput68 i_wb_we net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_116_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05607__A1 stack\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05607__B2 stack\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput79 rambus_wb_dat_i[10] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10529_ _00121_ clknet_leaf_113_clock mem.mem_dff.code_mem\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09349__A2 _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10054__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06032__A1 _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08309__B1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07740_ _02164_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08459__I _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__I mem.mem_dff.code_mem\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07671_ mem.mem_dff.code_mem\[31\]\[0\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _04377_ _04365_ _04383_ _04385_ _04375_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06622_ _02064_ _02118_ _02130_ _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06553_ mem.mem_dff.code_mem\[1\]\[1\] _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09341_ _03242_ _04319_ _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_169_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05504_ _01040_ _01047_ _01052_ _01053_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06484_ _02014_ _02015_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09272_ net256 _04256_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08223_ mem.mem_dff.data_mem\[0\]\[2\] _03318_ _03319_ _03416_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05435_ _00984_ _00985_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_194_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__A1 _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08154_ _02097_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05366_ _00918_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ _02512_ _02502_ _02513_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08085_ net75 _03273_ _03274_ net126 _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05297_ _00850_ _00776_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ mem.mem_dff.code_mem\[13\]\[5\] _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06271__A1 _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input40_I i_wb_addr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08987_ _03973_ _04043_ _04044_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07938_ _03154_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09512__A2 _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10542__CLK clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output127_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ _03109_ _03103_ _03110_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ _04544_ cycles_per_ms\[11\] _04567_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10880_ _00472_ clknet_leaf_148_clock stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09539_ delay_cycles\[23\] _04498_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__A2 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06617__I mem.mem_dff.code_mem\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10692__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10139__I _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09928__I _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09579__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11048__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09043__A4 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10314_ _03882_ _05117_ _05127_ _05128_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06352__I _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__B1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10245_ _04218_ _05074_ _05078_ stack\[14\]\[1\] _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05860__I1 stack\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09200__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ net169 _05023_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05999__S1 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06301__B _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07911__I mem.mem_dff.data_mem\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_170_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07817__A2 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09019__A1 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09838__I _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05220_ net136 _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08778__B1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_1_0_clock clknet_0_clock clknet_2_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10415__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06253__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09990__A2 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ net151 _03974_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09890_ _04799_ _04800_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_95_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05807__S _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09742__A2 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08545__A3 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _03932_ _03933_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10565__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__B1 _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ _03879_ _03871_ _03880_ _03881_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05984_ _01521_ _01527_ _00852_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05764__B1 _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ mem.mem_dff.data_mem\[0\]\[2\] _02992_ _02982_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07654_ _02928_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08917__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05516__B1 _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07821__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06605_ _02116_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09258__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07585_ _02877_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08138__B _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09324_ _04270_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06536_ _02058_ _02049_ _02061_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _04225_ _04235_ _04242_ stack\[22\]\[4\] _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06467_ _01995_ _02001_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ mem.mem_dff.code_mem\[11\]\[2\] _02383_ _02815_ mem.mem_dff.code_mem\[26\]\[2\]
+ _03399_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05295__A2 _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input88_I rambus_wb_dat_i[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05418_ stack\[19\]\[3\] stack\[16\]\[3\] stack\[17\]\[3\] stack\[18\]\[3\] _00968_
+ _00969_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09186_ _04190_ _04194_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06398_ _01425_ _01447_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_162_clock clknet_4_3_0_clock clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ _03317_ _03332_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05349_ _00883_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06244__A1 _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06172__I _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08068_ net115 _03250_ _03268_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__A1 _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07019_ _02351_ _02446_ _02437_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_177_clock clknet_4_4_0_clock clknet_leaf_177_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10030_ delay_counter\[4\] _04901_ _04882_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09733__A2 _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07744__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_3_0_clock clknet_3_1_0_clock clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_100_clock clknet_4_13_0_clock clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09497__A1 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10932_ _00524_ clknet_leaf_191_clock stack\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _00455_ clknet_leaf_144_clock stack\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09249__A1 _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_115_clock clknet_4_12_0_clock clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _00386_ clknet_leaf_170_clock stack\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10438__CLK clknet_leaf_75_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05905__S1 _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06483__A1 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06082__I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_117_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10319__B1 _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09185__B1 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _01963_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08932__B1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _05012_ _05014_ _05010_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _02370_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06257__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08999__B1 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09040_ _04038_ _04082_ _04083_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06252_ stack\[2\]\[1\] _01718_ _01793_ _01759_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08472__I _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05203_ mem.addr\[1\] _00757_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01724_ _01725_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06226__A1 _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10022__A2 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_94_clock clknet_4_13_0_clock clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06777__A2 _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _04798_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09715__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _04784_ _04789_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05764__C _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _03917_ _03921_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05336__I _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _01762_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05967_ _01390_ _01509_ _01510_ _01394_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09479__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ _02981_ _02973_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_clock clknet_4_10_0_clock clknet_leaf_32_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _03789_ _03809_ _03812_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05898_ _00790_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06001__I1 stack\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ _02928_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07568_ _02875_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09100__B1 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ net100 _02289_ _00760_ net96 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06519_ _02043_ _02029_ _02047_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_47_clock clknet_4_9_0_clock clknet_leaf_47_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _02737_ _02819_ _02810_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ _04137_ _04229_ _04208_ _04112_ _04231_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_output194_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10730__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08206__A2 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09403__A1 _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ _04131_ _04161_ _04178_ stack\[1\]\[5\] _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11200_ net110 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06217__B2 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09954__A2 _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07965__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11131_ _00723_ clknet_leaf_173_clock stack\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10880__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11062_ _00654_ clknet_leaf_21_clock delay_cycles\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08914__B1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _04881_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05246__I _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06940__A2 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__B _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10915_ _00507_ clknet_leaf_188_clock stack\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09890__A1 _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08693__A2 _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _00438_ clknet_leaf_161_clock stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ _00369_ clknet_leaf_53_clock net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06456__A1 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__I mem.mem_dff.code_mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10252__A2 _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06456__B2 stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06208__A1 _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10004__A2 _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06759__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__A1 _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06540__I _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ mem.mem_dff.code_mem\[9\]\[2\] _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09851__I _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05821_ stack\[20\]\[7\] stack\[21\]\[7\] _01360_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08540_ _01964_ _03693_ _03695_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05752_ stack\[18\]\[2\] stack\[19\]\[2\] stack\[16\]\[2\] stack\[17\]\[2\] _00792_
+ _00884_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08467__I _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _03636_ _03637_ _01692_ _03640_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05683_ _01190_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09881__A1 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__A2 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06695__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ _02761_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05498__A2 stack\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07353_ _02626_ _02705_ _02697_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10753__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07239__A3 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06304_ _00981_ _01841_ _01843_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10243__A2 _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ mem.mem_dff.code_mem\[20\]\[1\] _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08987__A3 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _04071_ _04069_ _04072_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06235_ _01740_ _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11109__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08930__I _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06166_ _01606_ _01707_ _01647_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_219_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06097_ _01618_ _01640_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_160_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06450__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09925_ delay_cycles\[6\] _04824_ _04820_ _04827_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09856_ _04565_ _04767_ _04775_ net44 _03262_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08372__B2 mem.mem_dff.data_mem\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _03794_ _03892_ _03907_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _04412_ _04666_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06383__B1 _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06999_ _02427_ _02428_ _02430_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _01989_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08124__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output207_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _03736_ _03797_ _03799_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09872__B2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10700_ _00292_ clknet_leaf_66_clock mem.mem_dff.data_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05489__A2 _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10631_ _00223_ clknet_leaf_101_clock mem.mem_dff.code_mem\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10562_ _00154_ clknet_leaf_80_clock mem.mem_dff.code_mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06625__I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09001__I _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06989__A2 _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10493_ _00085_ clknet_leaf_120_clock mem.mem_dff.code_mem\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05949__B1 _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05413__A2 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11114_ _00706_ clknet_leaf_192_clock stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11045_ _00637_ clknet_leaf_26_clock delay_cycles\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10626__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08363__A1 mem.mem_dff.code_mem\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08363__B2 mem.mem_dff.code_mem\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_0_0_clock clknet_2_0_0_clock clknet_3_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05972__I0 stack\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10776__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09863__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A2 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09863__B2 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06677__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10829_ _00421_ clknet_leaf_157_clock stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06429__A1 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07140__B _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09091__A2 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ stack\[10\]\[1\] stack\[11\]\[1\] _01472_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08750__I _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07366__I _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05404__A2 _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06270__I _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07971_ mem.mem_dff.data_mem\[7\]\[7\] _03179_ _03183_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09710_ _04276_ _04297_ _04311_ _04344_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_06922_ mem.mem_dff.code_mem\[10\]\[5\] _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09146__A3 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xspell_269 rambus_wb_addr_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09641_ _04600_ _04596_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06853_ _02128_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10161__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05804_ _00832_ stack\[10\]\[0\] _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ delay_cycles\[12\] _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06784_ _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _03650_ _03677_ _03682_ stack\[29\]\[1\] _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05735_ _01278_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09854__A1 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09854__B2 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input105_I rambus_wb_dat_i[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08454_ _01631_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05666_ _01205_ _01209_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_212_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _02745_ _02746_ _02748_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08409__A2 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _03572_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09606__A1 _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05597_ _01144_ stack\[8\]\[7\] stack\[9\]\[7\] _01131_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07336_ mem.mem_dff.code_mem\[21\]\[6\] _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10216__A2 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05891__A2 _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05489__C _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _02522_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04011_ _04043_ _04057_ stack\[25\]\[4\] _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06218_ _01183_ _01642_ _01760_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05643__A2 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07198_ _02533_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11081__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06149_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07276__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10649__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08593__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06180__I _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output157_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09908_ delay_cycles\[2\] _04811_ _04808_ _04814_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09839_ _04766_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10152__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__C _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09845__A1 _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10614_ _00206_ clknet_leaf_107_clock mem.mem_dff.code_mem\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06355__I _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _00137_ clknet_leaf_96_clock mem.mem_dff.code_mem\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__I stack\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10476_ _00068_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08033__B1 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10391__A1 _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 mem.mem_dff.code_mem\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__B2 mem.mem_dff.code_mem\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _00620_ clknet_leaf_19_clock cycles_per_ms\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06347__B1 _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08887__A2 _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A1 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05570__A1 _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05520_ _01061_ _01069_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07311__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05451_ _00933_ _01001_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08170_ _02172_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05382_ _00933_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_220_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _02063_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07075__A1 _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08811__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ _02350_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06822__A1 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput112 net112 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06003_ _01272_ _01545_ _01546_ _01390_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput123 net123 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput134 net134 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput145 net145 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput156 net156 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput167 net167 o_wb_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput178 net178 o_wb_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput189 net189 rambus_wb_addr_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10382__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10941__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07954_ _02984_ _03171_ _03173_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08327__B2 mem.mem_dff.code_mem\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _02354_ _02349_ _02355_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07885_ _03122_ _03117_ _03113_ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10134__A1 _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08878__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__B2 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09624_ delay_cycles\[0\] _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06836_ _02300_ _02295_ _02301_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09555_ _04509_ _04493_ delay_cycles\[17\] _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06767_ _02121_ _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09827__A1 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08506_ _03628_ _01707_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_169_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05718_ stack\[2\]\[2\] stack\[3\]\[2\] stack\[0\]\[2\] stack\[1\]\[2\] _01261_ _00902_
+ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _04440_ _03628_ _04451_ _04453_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06698_ _02161_ _02187_ _02183_ _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08437_ _02051_ _03609_ _03611_ _03612_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05649_ net258 net158 _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08368_ _03553_ _03554_ _03555_ _03556_ _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _02626_ _02679_ _02672_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__B1 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08299_ mem.mem_dff.code_mem\[10\]\[5\] _03343_ _03344_ mem.mem_dff.code_mem\[24\]\[5\]
+ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08802__A2 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08390__I _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10330_ _05140_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _01676_ _03701_ _03994_ _03945_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_105_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10192_ net174 _05035_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10373__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10125__A1 _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__B2 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__A4 _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__I _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__A1 _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08565__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10814__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput14 i_la_data[6] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07057__A1 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput25 i_wb_addr[16] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 i_wb_addr[4] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput47 i_wb_data[13] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput58 i_wb_data[23] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05607__A2 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput69 io_in[0] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06813__I _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _00120_ clknet_leaf_113_clock mem.mem_dff.code_mem\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _00051_ clknet_leaf_72_clock mem.mem_dff.code_mem\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05429__I _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10364__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05791__A1 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _02951_ _02942_ _02954_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06621_ _02129_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A1 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05543__A1 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ mem.io_data_out\[4\] _04320_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06552_ _02068_ _02073_ _02075_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05503_ _00974_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09271_ _04252_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_91_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06483_ _00764_ _01175_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08222_ _03413_ _03414_ _03415_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10494__CLK clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05434_ _00968_ stack\[4\]\[4\] stack\[5\]\[4\] _00928_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09037__A2 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ mem.mem_dff.code_mem\[11\]\[1\] _02383_ _02815_ mem.mem_dff.code_mem\[26\]\[1\]
+ _03347_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05365_ _00917_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07104_ _02494_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _03281_ _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05296_ net140 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07035_ _02455_ _02456_ _02458_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06271__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10355__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _03679_ _03939_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input33_I i_wb_addr[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07937_ _02998_ _03155_ _03161_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ _03079_ _03104_ _03095_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_217_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06819_ net187 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09607_ _04545_ _04533_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07799_ _03053_ _03046_ _03055_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09538_ delay_cycles\[22\] _04497_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08385__I _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__B _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10837__CLK clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09469_ _04338_ _01668_ _04360_ _04437_ _03625_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_185_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09028__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10987__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05958__B _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ stack\[27\]\[5\] _05112_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10155__I _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08539__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08539__B2 stack\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _03890_ _05072_ _05079_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10346__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09200__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10175_ _05024_ _05026_ _05022_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05773__A1 _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08172__C1 mem.mem_dff.code_mem\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_113_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09019__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08778__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08778__B2 stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05587__C _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06253__A2 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11142__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ net149 _03930_ _03928_ stack\[7\]\[5\] _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__B2 stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08771_ _03762_ _03864_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05983_ _01355_ _01523_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07722_ _02108_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ mem.mem_dff.code_mem\[30\]\[4\] _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09522__C _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05516__A1 stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05516__B2 _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06604_ net240 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07584_ mem.mem_dff.code_mem\[28\]\[4\] _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09258__A2 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05622__I _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ net103 _04304_ _02134_ net97 _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_209_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06535_ _02060_ _02052_ _02046_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04175_ _04234_ _04243_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06466_ mem.dff_data_ready _01996_ _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08205_ _03396_ _03397_ _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08218__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05417_ _00962_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06492__A2 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09185_ _04191_ _04192_ _04193_ _04167_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06397_ _01932_ _01933_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08136_ mem.mem_dff.data_mem\[0\]\[0\] _03318_ _03319_ _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05348_ _00900_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07441__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_3_0_clock_I clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06244__A2 _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ net72 _03252_ _03254_ net123 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05279_ stack\[19\]\[0\] stack\[16\]\[0\] stack\[17\]\[0\] stack\[18\]\[0\] _00821_
+ _00828_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09764__I _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07018_ _02444_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A2 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09194__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07744__A2 _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _04006_ _04028_ _04030_ stack\[0\]\[2\] _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _00523_ clknet_leaf_182_clock stack\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05507__A1 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _00454_ clknet_leaf_152_clock stack\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11015__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _00385_ clknet_leaf_169_clock stack\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09939__I _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09957__B1 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06363__I _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07432__A1 _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05294__I0 stack\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05908__S _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10319__A1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09185__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _05064_ _05054_ _05065_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09185__B2 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08932__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08932__B2 stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10158_ _04551_ _05008_ _05013_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10089_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07499__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05442__I _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08999__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06320_ _01023_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__B2 stack\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05357__S0 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09660__A2 _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06251_ _01792_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07369__I mem.mem_dff.code_mem\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05202_ _00760_ net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09948__B1 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06273__I _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ net8 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07423__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05818__S _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05434__B1 stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _04829_ _04839_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09872_ cycles_per_ms\[16\] _04785_ _04788_ net50 _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10682__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08923__A1 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _03918_ _03919_ _03920_ _03866_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08754_ _03863_ _03867_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05966_ stack\[14\]\[4\] stack\[15\]\[4\] _01369_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09479__A2 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07832__I mem.mem_dff.data_mem\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07705_ _02952_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11038__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08685_ _03654_ _03805_ _03803_ stack\[5\]\[3\] _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05897_ stack\[4\]\[6\] stack\[5\]\[6\] _00881_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08151__A2 _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07636_ _02874_ _02927_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06162__A1 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07567_ _02760_ _02813_ _02171_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09759__I _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _01196_ _04265_ _04287_ _04289_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06518_ _02045_ _02032_ _02046_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09100__B2 stack\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07498_ mem.mem_dff.code_mem\[26\]\[1\] _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ stack\[21\]\[7\] _04213_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06449_ _01984_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10261__A3 _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09168_ _03728_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output187_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ _03298_ _03305_ _03313_ _03314_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__06217__A2 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _01887_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11130_ _00722_ clknet_leaf_173_clock stack\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__I mem.mem_dff.code_mem\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05976__A1 _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05976__B2 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _00653_ clknet_leaf_21_clock delay_cycles\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05291__I3 stack\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05527__I _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08914__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04880_ _04886_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08914__B2 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09443__B _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10914_ _00506_ clknet_leaf_184_clock stack\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10845_ _00437_ clknet_leaf_161_clock stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05900__A1 _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05900__B2 _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _00368_ clknet_leaf_122_clock net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05339__S0 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10555__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06456__A2 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06026__C _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05967__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05967__B2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08905__A1 _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05719__A1 _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _00803_ _01361_ _01362_ _01363_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05881__B _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05751_ _01277_ _01294_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_161_clock clknet_4_6_0_clock clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _01711_ _03639_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06144__A1 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05682_ _01221_ _01225_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_208_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ _02760_ _02291_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ mem.mem_dff.code_mem\[22\]\[1\] _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_176_clock clknet_4_4_0_clock clknet_leaf_176_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06303_ _00981_ _01841_ _01842_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _02647_ _02652_ _02654_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09022_ _03996_ _03822_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06234_ _01771_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06165_ _01606_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_219_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05775__C _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06096_ _01639_ _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_114_clock clknet_4_12_0_clock clknet_leaf_114_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _04576_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09855_ _04778_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08806_ _03844_ _03893_ _03903_ stack\[6\]\[5\] _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10428__CLK clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _04724_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06998_ _02366_ _02429_ _02425_ _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07562__I _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_129_clock clknet_4_9_0_clock clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ _03846_ _03850_ _03852_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05949_ _01363_ _01491_ _01492_ _00844_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__A2 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ _03696_ _03773_ _03792_ stack\[4\]\[7\] _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06135__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__I _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09872__A2 _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10578__CLK clknet_leaf_89_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07619_ _02903_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _03740_ _03742_ _03744_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_148_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10219__B1 _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10630_ _00222_ clknet_leaf_102_clock mem.mem_dff.code_mem\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ _00153_ clknet_leaf_96_clock mem.mem_dff.code_mem\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08832__B1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _00084_ clknet_leaf_120_clock mem.mem_dff.code_mem\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05249__I0 stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05949__A1 _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05949__B2 _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _00705_ clknet_leaf_178_clock stack\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05413__A3 stack\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ _00636_ clknet_4_2_0_clock delay_cycles\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08363__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05972__I1 stack\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08115__A2 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09312__A1 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_clock clknet_4_13_0_clock clknet_leaf_93_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09863__A2 _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05921__S _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ _00420_ clknet_leaf_171_clock stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05720__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06429__A2 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__B1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10759_ _00351_ clknet_leaf_49_clock mem.dff_data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_31_clock clknet_4_10_0_clock clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08051__A1 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08051__B2 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06601__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07970_ _03167_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_214_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06921_ _02363_ _02364_ _02368_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_46_clock clknet_4_9_0_clock clknet_leaf_46_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xspell_259 o_wb_data[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06852_ mem.mem_dff.code_mem\[8\]\[7\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09640_ cycles_per_ms\[1\] _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08478__I _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05799__S0 _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05803_ stack\[11\]\[0\] _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09571_ delay_cycles\[15\] _04530_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06783_ _02169_ _02258_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10720__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08106__A2 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09303__A1 _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05963__I1 stack\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08522_ _01183_ _03671_ _03683_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_188_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05734_ _01274_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09854__A2 _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05831__S _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08453_ _03622_ _03623_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07865__A1 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05665_ _01189_ _01206_ _01208_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_212_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_161_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ _02717_ _02747_ _02743_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06726__I _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ _03571_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05596_ _01083_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09606__A2 _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__I _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _02692_ _02689_ _02693_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__B1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09082__A3 _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07266_ mem.mem_dff.code_mem\[19\]\[6\] _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08290__A1 _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__I _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09005_ _01860_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06217_ stack\[2\]\[0\] _01718_ _01758_ _01759_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07197_ mem.mem_dff.code_mem\[18\]\[0\] _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input63_I i_wb_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06148_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08593__A2 _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06079_ net256 _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_86_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ _04590_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_154_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08345__A2 _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08388__I _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _04766_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05403__I0 stack\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09769_ exec.memory_input\[4\] _04322_ _04715_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05540__I _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10613_ _00205_ clknet_leaf_106_clock mem.mem_dff.code_mem\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ _00136_ clknet_leaf_97_clock mem.mem_dff.code_mem\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08851__I _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10475_ _00067_ clknet_leaf_123_clock mem.mem_dff.code_mem\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08033__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08033__B2 stack\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A2 _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10743__CLK clknet_leaf_167_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11027_ _00619_ clknet_leaf_17_clock cycles_per_ms\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__B _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05715__I _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05570__A2 _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout250_I net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05450_ _00942_ stack\[20\]\[4\] stack\[21\]\[4\] _00962_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05381_ _00923_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ mem.mem_dff.code_mem\[15\]\[7\] _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _02470_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07377__I _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06002_ stack\[20\]\[1\] stack\[21\]\[1\] _01329_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput113 net113 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput124 net124 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput135 net135 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_108_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput146 net146 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput157 net157 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net168 o_wb_data[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput179 net179 o_wb_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A2 _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05826__S _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ mem.mem_dff.data_mem\[7\]\[0\] _03172_ _03168_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06904_ _02264_ _02352_ _02342_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07884_ _02059_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A1 _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05625__I mem.sram_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09623_ delay_cycles\[1\] _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08001__I _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06835_ _02235_ _02296_ _02283_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06766_ mem.mem_dff.code_mem\[6\]\[5\] _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09554_ cycles_per_ms\[17\] _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05717_ _00881_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08505_ _01991_ _03665_ _03667_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06697_ mem.mem_dff.code_mem\[4\]\[6\] _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09485_ _01064_ _04441_ _04452_ _04339_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07061__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08436_ _02009_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05648_ net129 _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08367_ mem.mem_dff.code_mem\[3\]\[7\] _03364_ _03365_ mem.mem_dff.code_mem\[4\]\[7\]
+ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05579_ _01102_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07318_ mem.mem_dff.code_mem\[21\]\[1\] _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10616__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A1 mem.mem_dff.code_mem\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08298_ mem.mem_dff.code_mem\[8\]\[5\] _02293_ _02701_ mem.mem_dff.code_mem\[22\]\[5\]
+ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07249_ _02625_ _02622_ _02627_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10260_ _04205_ _05086_ _05088_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10766__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _05036_ _05038_ _05034_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10373__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A2 _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06329__A1 _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05535__I _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08846__I _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__I _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 i_la_data[7] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput26 i_wb_addr[17] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput37 i_wb_addr[5] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 i_wb_data[14] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10061__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput59 i_wb_data[2] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _00119_ clknet_leaf_112_clock mem.mem_dff.code_mem\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10458_ _00050_ clknet_leaf_70_clock mem.mem_dff.code_mem\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__A2 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10389_ stack\[15\]\[3\] _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10364__A2 _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__A2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__A1 _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10116__A2 _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06620_ _02128_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08756__I _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07660__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09809__A2 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11071__CLK clknet_opt_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _02031_ _02074_ _02066_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05502_ _01009_ _01048_ _01050_ _01051_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10639__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _04250_ _04251_ _04252_ _04254_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_21_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ _01994_ _02013_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08221_ mem.mem_dff.data_mem\[4\]\[2\] _03101_ _03131_ mem.mem_dff.data_mem\[5\]\[2\]
+ _03381_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05433_ _00923_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _03342_ _03345_ _03346_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08245__A1 mem.mem_dff.code_mem\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__I _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05364_ _00916_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07103_ _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10052__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08083_ _03261_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09993__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05295_ _00819_ _00848_ _00807_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_3_3_0_clock_I clknet_2_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _02366_ _02457_ _02453_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10355__A2 _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ _03672_ _03993_ _03944_ _03675_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07936_ mem.mem_dff.data_mem\[6\]\[3\] _03156_ _03160_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input26_I i_wb_addr[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ mem.mem_dff.data_mem\[4\]\[2\] _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09606_ _04565_ _04563_ _04561_ cycles_per_ms\[9\] _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06818_ _02017_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07798_ _02968_ _03047_ _03054_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09537_ delay_cycles\[21\] delay_cycles\[20\] _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06749_ mem.mem_dff.code_mem\[6\]\[1\] _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09468_ _01696_ _04411_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10291__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08419_ net127 _03125_ _03591_ _03592_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_145_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ _04359_ _04365_ _04366_ _04373_ _04375_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_162_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10043__B2 _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__A1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06798__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06135__B _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ _03228_ _05109_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08539__A2 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _01758_ _05074_ _05078_ stack\[14\]\[0\] _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07745__I mem.mem_dff.data_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10174_ cycles_per_ms\[16\] _05020_ _05025_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05222__A1 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10171__I _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05265__I _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__A2 _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11094__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08172__B1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__C2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06722__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10120__B _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06096__I _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A1 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09019__A3 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08227__B2 mem.mem_dff.code_mem\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08778__A2 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06045__B _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08950__A2 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05982_ _01401_ _01524_ _01525_ _01272_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08770_ stack\[11\]\[4\] _03872_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05764__A2 _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ _02994_ _02991_ _02995_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_211_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06013__I0 stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_10_0_clock_I clknet_3_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10461__CLK clknet_leaf_72_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _02938_ _02929_ _02940_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05516__A2 _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07390__I _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06603_ _02099_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07583_ _02885_ _02878_ _02887_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06534_ _02059_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09322_ _00758_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10273__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04222_ _04236_ _04242_ stack\[22\]\[3\] _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06465_ _01999_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08204_ mem.mem_dff.code_mem\[12\]\[2\] _02414_ _02442_ mem.mem_dff.code_mem\[13\]\[2\]
+ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05416_ _00945_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09184_ _04187_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06396_ _01713_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09110__I _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _03322_ _03326_ _03330_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09966__A1 _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05347_ _00899_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ _03243_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05278_ stack\[23\]\[0\] stack\[20\]\[0\] stack\[21\]\[0\] stack\[22\]\[0\] _00832_
+ _00823_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07017_ _02444_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05452__A1 stack\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05452__B2 stack\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07992__A3 _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__A2 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09194__A2 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_7_0_clock_I clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08968_ _03952_ _04023_ _04032_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output132_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07919_ mem.mem_dff.data_mem\[5\]\[6\] _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08899_ _03975_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10930_ _00522_ clknet_leaf_182_clock stack\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05813__I _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _00453_ clknet_leaf_145_clock stack\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10954__CLK clknet_leaf_179_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08457__A1 _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10792_ _00384_ clknet_leaf_159_clock stack\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10264__A1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__I _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__A1 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09957__B2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09709__A1 _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05443__A1 stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05294__I1 stack\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08080__B _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09185__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10226_ _04227_ _05045_ _05062_ stack\[12\]\[5\] _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10157_ _04950_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08932__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A1 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05924__S _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10088_ _04955_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06819__I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05723__I _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10255__A1 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__S1 _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06250_ _01791_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05598__C _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05201_ _00759_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06181_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09865__I _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05434__A1 _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09940_ _04545_ _04835_ _04832_ _04838_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05434__B2 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07385__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10827__CLK clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _04774_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08923__A2 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _03914_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09814__B _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06934__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08753_ _03208_ _03864_ _03865_ _03866_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05965_ stack\[12\]\[4\] stack\[13\]\[4\] _01391_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ _02063_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05896_ _01313_ _01439_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08684_ _03787_ _03809_ _03811_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09105__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07635_ _02926_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08439__A1 _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _02531_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08944__I _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _04288_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10246__A1 _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09100__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06517_ _01999_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07497_ _02812_ _02817_ _02820_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I rambus_wb_dat_i[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06464__I _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _04133_ _04229_ _04230_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06448_ _01216_ _01820_ _01821_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10261__A4 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09167_ _04177_ _04171_ _04179_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06379_ _01890_ _01904_ _01809_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_175_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ mem.mem_dff.code_mem\[7\]\[0\] _02258_ _02469_ mem.mem_dff.code_mem\[14\]\[0\]
+ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ _04056_ _04115_ _04128_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05425__A1 _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08049_ _02291_ _03248_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05808__I stack\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11060_ _00652_ clknet_leaf_22_clock delay_cycles\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09167__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_156_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ delay_counter\[1\] _04647_ _04885_ _00876_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06925__A1 _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05744__S _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ _00505_ clknet_leaf_178_clock stack\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07350__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11132__CLK clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10844_ _00436_ clknet_leaf_189_clock stack\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08854__I _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _00367_ clknet_leaf_122_clock net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05339__S1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05967__A2 _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08366__B1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10209_ _05049_ _05052_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08905__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11189_ net237 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05719__A2 stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05750_ _01279_ _01293_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06549__I _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__A1 _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05681_ _01224_ _01194_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07341__A1 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _02022_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_211_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__B1 _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _02699_ _02703_ _02706_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09094__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06302_ _01236_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ _02591_ _02653_ _02645_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06284__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09021_ _03780_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06233_ _00875_ _01772_ _01773_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09809__B _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06164_ _01620_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10400__A1 _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06095_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05958__A2 stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06080__A1 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09923_ _04816_ _04826_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11005__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09854_ _04559_ _04767_ _04775_ net66 _03262_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__I _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _03791_ _03901_ _03906_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09785_ _04724_ _04726_ _04727_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08109__B1 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06997_ _02416_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06383__A2 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ _03851_ _03831_ _03840_ stack\[8\]\[6\] _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11155__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05948_ stack\[26\]\[4\] stack\[27\]\[4\] _01369_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05591__B1 stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ _03732_ _03797_ _03798_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05879_ _01408_ _01415_ _01421_ _01422_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07618_ mem.mem_dff.code_mem\[29\]\[4\] _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _01618_ _03743_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07549_ _02847_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09085__A1 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_82_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06194__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10560_ _00152_ clknet_leaf_96_clock mem.mem_dff.code_mem\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08832__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08832__B2 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _04218_ _04215_ _04213_ stack\[21\]\[1\] _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ _00083_ clknet_leaf_120_clock mem.mem_dff.code_mem\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05739__S _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07399__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05538__I _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11112_ _00704_ clknet_leaf_178_clock stack\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11043_ _00635_ clknet_leaf_26_clock delay_cycles\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05257__S0 _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09560__A2 _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05421__I1 stack\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10522__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06126__A2 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08584__I _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09076__A1 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ _00419_ clknet_leaf_171_clock stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10758_ _00350_ clknet_leaf_47_clock mem.dff_data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08823__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08823__B2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10689_ _00281_ clknet_leaf_67_clock mem.mem_dff.data_mem\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07928__I _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09379__A2 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11028__CLK clknet_leaf_19_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06920_ _02366_ _02367_ _02361_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06851_ _02311_ _02306_ _02312_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05799__S1 _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05802_ stack\[8\]\[0\] stack\[9\]\[0\] _00822_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _04487_ _04488_ _04492_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06279__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06782_ _02257_ _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__A2 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ _03633_ _03677_ _03682_ stack\[29\]\[0\] _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05733_ _01260_ _01262_ _01276_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07612__B _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_104_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _01769_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05664_ _01190_ _01207_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _02732_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08383_ _02813_ _02986_ _03247_ _03570_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__09067__A1 stack\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05595_ _01129_ _01139_ _01142_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07334_ _02608_ _02690_ _02686_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08814__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08814__B2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05628__A1 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__A4 _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ _02638_ _02635_ _02639_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_192_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07838__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09004_ _04056_ _04052_ _04058_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06216_ _01714_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07196_ _02582_ _02575_ _02584_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ _01686_ _01688_ _01689_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input56_I i_wb_data[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06078_ net110 _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05800__A1 _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ _04799_ _04813_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09837_ _01694_ _04362_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10545__CLK clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _04717_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _03787_ _03826_ _03838_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _04658_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06108__A2 _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__B1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10695__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07856__A2 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09058__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10612_ _00204_ clknet_leaf_106_clock mem.mem_dff.code_mem\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08805__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05619__A1 _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _00135_ clknet_leaf_97_clock mem.mem_dff.code_mem\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07748__I _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10474_ _00066_ clknet_leaf_57_clock mem.mem_dff.code_mem\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_160_clock clknet_4_6_0_clock clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09230__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__A2 _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05268__I _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08579__I _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_175_clock clknet_4_4_0_clock clknet_leaf_175_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11026_ _00618_ clknet_leaf_17_clock cycles_per_ms\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06099__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05555__B1 stack\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06827__I _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07432__B _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__I _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_113_clock clknet_4_12_0_clock clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05380_ _00931_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_3_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10418__CLK clknet_leaf_39_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07050_ _02411_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_clock clknet_4_9_0_clock clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06001_ stack\[22\]\[1\] stack\[23\]\[1\] _00791_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput114 net114 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput125 net125 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_126_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput136 net136 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput158 net158 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10568__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput169 net169 o_wb_data[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_30_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07783__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07952_ _03170_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05794__B1 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__I mem.mem_dff.code_mem\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06903_ mem.mem_dff.code_mem\[10\]\[1\] _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_214_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ mem.mem_dff.data_mem\[4\]\[6\] _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06338__A2 _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09622_ _04574_ _04489_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06834_ mem.mem_dff.code_mem\[8\]\[2\] _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05546__B1 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09553_ _04507_ _04508_ _04511_ _04512_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06765_ _02240_ _02241_ _02244_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09288__A1 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input110_I reset vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08504_ net152 _03646_ _03657_ stack\[19\]\[7\] _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05716_ _01259_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09484_ _04442_ _01769_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06696_ _02189_ _02186_ _02190_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05641__I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08435_ net116 _03610_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05647_ _01190_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08366_ mem.mem_dff.code_mem\[19\]\[7\] _03366_ _03359_ mem.mem_dff.code_mem\[21\]\[7\]
+ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08248__C1 mem.mem_dff.code_mem\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__I _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05578_ _00950_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07317_ _02674_ _02678_ _02680_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _03485_ _03486_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08263__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _02626_ _02623_ _02615_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02557_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10358__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06026__A1 _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_92_clock clknet_4_13_0_clock clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10190_ cycles_per_ms\[20\] _05032_ _05037_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08971__B1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05816__I _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__A1 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06329__A2 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09451__C _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_30_clock clknet_4_11_0_clock clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10169__I _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_clock clknet_4_9_0_clock clknet_leaf_45_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08254__A2 _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 i_la_wb_disable net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 i_wb_addr[18] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07478__I mem.mem_dff.code_mem\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput38 i_wb_addr[6] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06265__A1 _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _00118_ clknet_leaf_111_clock mem.mem_dff.code_mem\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput49 i_wb_data[15] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__10061__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10710__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10457_ _00049_ clknet_leaf_70_clock mem.mem_dff.code_mem\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A2 _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10388_ _05179_ _05171_ _05180_ _05181_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05776__B1 _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10860__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__A2 _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07517__A1 _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11009_ _00601_ clknet_leaf_46_clock mem.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06740__A2 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07162__B _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06550_ _02072_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05461__I _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05501_ _00937_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06481_ net253 _01996_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08493__A2 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ mem.mem_dff.data_mem\[1\]\[2\] _03377_ _03378_ mem.mem_dff.data_mem\[3\]\[2\]
+ mem.mem_dff.data_mem\[7\]\[2\] _03379_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05432_ _00983_ net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ mem.mem_dff.code_mem\[12\]\[1\] _02414_ _02442_ mem.mem_dff.code_mem\[13\]\[1\]
+ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05363_ _00898_ _00915_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08245__A2 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__A3 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ _02044_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08082_ _03263_ _03280_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05294_ stack\[23\]\[1\] stack\[20\]\[1\] stack\[21\]\[1\] stack\[22\]\[1\] _00822_
+ _00847_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07033_ _02444_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05837__S _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_7_0_clock_I clknet_2_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08984_ _03936_ _04039_ _04042_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05636__I _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07935_ _03126_ _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08012__I _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _03106_ _03103_ _03108_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ cycles_per_ms\[10\] _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06817_ mem.mem_dff.code_mem\[8\]\[0\] _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input19_I i_wb_addr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ _03010_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ delay_cycles\[19\] _04485_ _04495_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06748_ _02223_ _02228_ _02231_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05790__I0 stack\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _04431_ _04384_ _04435_ _04436_ _04401_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06679_ mem.mem_dff.code_mem\[4\]\[1\] _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ net127 _03588_ _03589_ _03125_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__A2 _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _04374_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ mem.dff_data_out\[6\] _03538_ _03483_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__A2 _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09984__A2 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10311_ _03879_ _05117_ _05125_ _05126_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06930__I mem.mem_dff.code_mem\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _05077_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07747__A1 _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _04950_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05222__A2 _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_5_0_clock clknet_4_11_0_clock clknet_opt_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08857__I _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08172__A1 mem.mem_dff.code_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09688__I _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09019__A4 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10509_ _00101_ clknet_leaf_110_clock mem.mem_dff.code_mem\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__B1 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06410__A1 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05844__S0 _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05981_ stack\[22\]\[5\] stack\[23\]\[5\] _01403_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07720_ mem.mem_dff.data_mem\[0\]\[1\] _02992_ _02982_ _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10606__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07671__I mem.mem_dff.code_mem\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06013__I1 stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ _02857_ _02931_ _02939_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06602_ mem.mem_dff.code_mem\[2\]\[4\] _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07582_ _02857_ _02879_ _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_207_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09112__B1 _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09321_ _03622_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06533_ net235 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_14_0_clock_I clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10756__CLK clknet_leaf_48_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09663__A1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _04237_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10273__A2 _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08203_ mem.mem_dff.code_mem\[25\]\[2\] _03340_ _03341_ mem.mem_dff.code_mem\[27\]\[2\]
+ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05415_ stack\[23\]\[3\] _00960_ _00961_ _00966_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_147_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09415__A1 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ _04186_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06395_ _01926_ _01931_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ mem.mem_dff.data_mem\[2\]\[0\] _03327_ _03329_ mem.mem_dff.data_mem\[6\]\[0\]
+ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05346_ _00785_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08007__I _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08065_ _03263_ _03266_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05277_ _00827_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_190_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07016_ _02411_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05452__A2 _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09718__A2 _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05794__C _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05366__I _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ _04004_ _04028_ _04030_ stack\[0\]\[1\] _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07918_ _03147_ _03144_ _03148_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08898_ _03952_ _03970_ _03978_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07581__I _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output125_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07849_ mem.mem_dff.data_mem\[3\]\[7\] _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10860_ _00452_ clknet_leaf_0_clock stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09103__B1 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09654__A1 _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_152_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10791_ _00383_ clknet_leaf_135_clock stack\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08457__A2 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05515__I0 stack\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__A2 _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09957__A2 _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__A2 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05818__I1 stack\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__I mem.mem_dff.data_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05294__I2 stack\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10225_ _03728_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10629__CLK clknet_leaf_102_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A1 _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_77_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10156_ net164 _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ net68 _01627_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07491__I _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10779__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A2 _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10989_ _00581_ clknet_leaf_40_clock mem.sram_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06459__A1 _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10255__A2 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05879__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__C _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06056__B _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05200_ mem.addr\[1\] mem.addr\[0\] _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05682__A2 _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _01625_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05434__A2 stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11188__I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09870_ _04784_ _04787_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08821_ _03913_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _00842_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05964_ _01409_ _01506_ _01507_ _01414_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07703_ mem.mem_dff.code_mem\[31\]\[7\] _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _03652_ _03805_ _03803_ stack\[5\]\[2\] _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09884__A1 _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05895_ stack\[2\]\[6\] stack\[3\]\[6\] stack\[0\]\[6\] stack\[1\]\[6\] _01438_ _00828_
+ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06698__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ _02787_ _02440_ _02224_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05745__I0 stack\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ mem.mem_dff.code_mem\[28\]\[0\] _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09304_ _02003_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07350__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06516_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10246__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06745__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07496_ _02818_ _02819_ _02810_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04135_ _04211_ _04223_ stack\[21\]\[6\] _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06447_ _01770_ _01972_ _01973_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input86_I rambus_wb_dat_i[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ _04129_ _04161_ _04178_ stack\[1\]\[4\] _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08960__I _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06378_ _01074_ _01811_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11084__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ mem.mem_dff.code_mem\[16\]\[0\] _02536_ _03307_ _03312_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_163_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05329_ _00881_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09097_ _04126_ _04117_ _04127_ stack\[24\]\[3\] _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06622__A1 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05425__A2 _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10010_ _04879_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10182__A1 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06386__B1 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _04870_ _01968_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09875__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ _00504_ clknet_leaf_178_clock stack\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10843_ _00435_ clknet_leaf_190_clock stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05361__A1 _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10774_ _00366_ clknet_leaf_53_clock net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__I _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10451__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__B _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09563__B1 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10208_ _04191_ _05050_ _05051_ _04167_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11188_ net241 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10139_ _04998_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05975__I0 stack\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05680_ _01223_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A1 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09618__B2 _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06565__I _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07170__B _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ _02704_ _02705_ _02697_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09094__A2 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ _00841_ _00875_ _00917_ _01840_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07281_ _02651_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09876__I _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _04069_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06232_ _00840_ _00875_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08780__I _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06163_ _01130_ _01705_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07396__I mem.mem_dff.code_mem\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10400__A2 _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06006__S _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _01621_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10944__CLK clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09922_ delay_cycles\[5\] _04824_ _04820_ _04825_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09853_ _04777_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10164__A1 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _03842_ _03893_ _03903_ stack\[6\]\[4\] _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09784_ _00764_ _04724_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06996_ _02416_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05966__I0 stack\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08735_ _03237_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08020__I _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05947_ stack\[24\]\[4\] stack\[25\]\[4\] _01391_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05591__A1 _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05591__B2 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__I0 stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08666_ _03694_ _03773_ _03792_ stack\[4\]\[6\] _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05878_ _01306_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07617_ _02911_ _02904_ _02913_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05343__A1 _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08597_ _03644_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10219__A2 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07548_ mem.mem_dff.code_mem\[27\]\[4\] _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06475__I _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09085__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07096__A1 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07479_ _02721_ _02803_ _02799_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08832__A2 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10474__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _01792_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _00082_ clknet_leaf_118_clock mem.mem_dff.code_mem\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _04161_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05249__I2 stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11111_ _00703_ clknet_leaf_151_clock stack\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__A1 _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11042_ _00634_ clknet_leaf_17_clock delay_cycles\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05257__S1 _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05554__I _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05421__I2 stack\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09848__A1 _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08086__B _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06385__I _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10826_ _00418_ clknet_leaf_169_clock stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10817__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10757_ _00349_ clknet_leaf_47_clock mem.dff_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08823__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10688_ _00280_ clknet_leaf_61_clock mem.mem_dff.data_mem\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10967__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__A1 stack\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08339__A1 _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__A2 _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06850_ _02279_ _02307_ _02303_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05948__I0 stack\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05464__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05801_ _01267_ _01340_ _01341_ _01342_ _01344_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06781_ _02025_ _02256_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05732_ _01263_ _01268_ _01269_ _01273_ _01275_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _03621_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05663_ _01192_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ _02732_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10497__CLK clknet_leaf_117_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06295__I _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08382_ net253 _00763_ _01177_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09067__A2 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05594_ stack\[14\]\[7\] _01140_ _01141_ stack\[15\]\[7\] _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07333_ mem.mem_dff.code_mem\[21\]\[5\] _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07078__A1 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08275__B1 _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ _02608_ _02636_ _02632_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09003_ _04008_ _04048_ _04057_ stack\[25\]\[3\] _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06215_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07195_ _02527_ _02576_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05639__I _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08015__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06146_ _01647_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _01603_ _01620_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07854__I _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09905_ _04583_ _04811_ _04808_ _04812_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input49_I i_wb_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__A2 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07075__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09836_ _04312_ _04758_ _04765_ _04761_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05939__I0 stack\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05374__I _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05403__I2 stack\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06979_ _02414_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09767_ exec.memory_input\[3\] _04311_ _04715_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ _03837_ _03830_ _03833_ stack\[8\]\[2\] _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04656_ _04657_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08502__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08502__B2 stack\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output205_I net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08649_ _03650_ _03779_ _03783_ stack\[4\]\[1\] _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09058__A2 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09302__I0 mem.io_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _00203_ clknet_leaf_107_clock mem.mem_dff.code_mem\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08805__A2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _00134_ clknet_leaf_97_clock mem.mem_dff.code_mem\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09449__C _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__B1 _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06292__A2 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10473_ _00065_ clknet_leaf_58_clock mem.mem_dff.code_mem\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09230__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _00617_ clknet_leaf_15_clock cycles_per_ms\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05284__I _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05555__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05555__B2 _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08595__I _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09049__A2 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _00401_ clknet_leaf_167_clock stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__I _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06843__I _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08009__B1 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11145__CLK clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__B _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05459__I _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06000_ _01313_ _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput115 net115 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_177_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10367__A1 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput126 net126 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput137 net137 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput148 net148 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_217_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput159 net258 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07783__A2 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ _03170_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10119__A1 _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11196__I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06902_ _02344_ _02349_ _02353_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07882_ _03119_ _03116_ _03120_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06833_ _02298_ _02295_ _02299_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09621_ cycles_per_ms\[5\] _04580_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05546__A1 _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05546__B2 stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09552_ cycles_per_ms\[19\] _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06764_ _02242_ _02243_ _02238_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08503_ _01964_ _03665_ _03666_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05715_ _01258_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09483_ _04402_ _04450_ _04414_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06695_ _02122_ _02187_ _02183_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _03601_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input103_I rambus_wb_dat_i[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05646_ net130 _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08365_ mem.mem_dff.code_mem\[2\]\[7\] _03349_ _03350_ mem.mem_dff.code_mem\[18\]\[7\]
+ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08248__B1 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08248__C2 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05577_ _01125_ net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07849__I mem.mem_dff.data_mem\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07316_ _02591_ _02679_ _02672_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06753__I _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ mem.mem_dff.code_mem\[23\]\[5\] _03391_ _03392_ mem.mem_dff.code_mem\[31\]\[5\]
+ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ _02505_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07471__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05369__I _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ mem.mem_dff.code_mem\[17\]\[3\] _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10358__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10512__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06129_ _01126_ _01670_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08971__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08971__B2 stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output155_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08723__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06329__A3 _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09771__I0 exec.memory_input\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09819_ net157 _04740_ _04741_ _04753_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_189_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05537__A1 _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09304__I _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0_clock clknet_4_0_0_clock clknet_opt_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_168_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08254__A3 _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09451__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 i_la_write net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput28 i_wb_addr[19] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_204_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 i_wb_addr[7] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10185__I _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _00117_ clknet_leaf_110_clock mem.mem_dff.code_mem\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10456_ _00048_ clknet_leaf_70_clock mem.mem_dff.code_mem\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10349__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10387_ _04100_ _05174_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07494__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_147_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09506__A3 _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11008_ _00600_ clknet_leaf_127_clock mem.mem_dff.memory_type_data vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06838__I _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__I _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05742__I _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05500_ stack\[30\]\[5\] _01049_ _00960_ stack\[31\]\[5\] _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06480_ mem.mem_dff.code_mem\[0\]\[0\] _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05431_ _00982_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05700__A1 _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ mem.mem_dff.code_mem\[10\]\[1\] _03343_ _03344_ mem.mem_dff.code_mem\[24\]\[1\]
+ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09978__B1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05362_ _00781_ _00909_ _00914_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_174_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09442__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ mem.mem_dff.code_mem\[15\]\[3\] _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08081_ mem.io_data_out\[5\] _03267_ _03271_ _03279_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05293_ _00802_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07032_ _02444_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10685__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__A1 stack\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06014__S _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05767__A1 _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08983_ _03937_ _04021_ _04035_ stack\[0\]\[7\] _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05311__S0 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07934_ _02996_ _03155_ _03159_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ _03107_ _03104_ _03095_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ cycles_per_ms\[10\] _04563_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07353__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06816_ _02281_ _02273_ _02284_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07796_ mem.mem_dff.data_mem\[2\]\[3\] _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05652__I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06747_ _02229_ _02230_ _02221_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09535_ _04494_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05790__I1 stack\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _04357_ _04399_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06678_ _02168_ _02175_ _02177_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _03594_ _03597_ _03598_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05629_ mem.mem_dff.memory_type_data _01175_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ _01644_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ _03532_ _03537_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08279_ mem.mem_dff.code_mem\[7\]\[4\] _03428_ _03432_ mem.mem_dff.code_mem\[14\]\[4\]
+ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _03762_ _05114_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05455__B1 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09197__A1 _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_189_clock clknet_4_1_0_clock clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10241_ _05075_ _05073_ _05076_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07747__A2 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ net168 _05023_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_112_clock clknet_4_12_0_clock clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08172__A2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10408__CLK clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_127_clock clknet_4_9_0_clock clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08873__I _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_73_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__I _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05511__B _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__I _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _00100_ clknet_leaf_108_clock mem.mem_dff.code_mem\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ _00031_ clknet_leaf_68_clock mem.mem_dff.code_mem\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__A1 _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08935__B2 stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05749__A1 _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05980_ stack\[20\]\[5\] stack\[21\]\[5\] _00791_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05844__S1 _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__I _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__B _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _02897_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06568__I mem.mem_dff.code_mem\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06174__A1 _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06601_ _02111_ _02100_ _02113_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07581_ _02841_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05405__C _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09320_ _01207_ _04265_ _04302_ _04289_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09112__A1 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ mem.mem_dff.code_mem\[0\]\[6\] _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10258__B1 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08783__I _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_clock clknet_4_15_0_clock clknet_leaf_91_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_179_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _04173_ _04234_ _04241_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07674__A1 _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ _01997_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08871__B1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08202_ mem.mem_dff.code_mem\[10\]\[2\] _02347_ _02762_ mem.mem_dff.code_mem\[24\]\[2\]
+ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05414_ _00934_ _00964_ _00965_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09182_ _03207_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06009__S _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06394_ _01930_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08133_ _03328_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07426__A1 _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05345_ _00879_ _00888_ _00897_ _00854_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05437__B1 stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05848__S _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ mem.io_data_out\[2\] _03244_ _03246_ _03265_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05276_ _00819_ _00824_ _00830_ _00816_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_190_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07015_ _02442_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08926__A1 stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__I _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08966_ _03819_ _04023_ _04031_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08958__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input31_I i_wb_addr[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07917_ _03090_ _03145_ _03141_ _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_44_clock clknet_4_9_0_clock clknet_leaf_44_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08897_ _03835_ _03972_ _03976_ stack\[10\]\[1\] _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08179__B _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09351__A1 _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07083__B _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07848_ _03092_ _03085_ _03093_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05382__I _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output118_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07779_ _02981_ _03032_ _03039_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09789__I _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09103__B2 stack\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _04252_ _04478_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_59_clock clknet_4_14_0_clock clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10790_ _00382_ clknet_leaf_135_clock stack\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ _04369_ _04419_ _04420_ _04382_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10850__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07102__I _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05279__I0 stack\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08090__A1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05979__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__C _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05294__I3 stack\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _05061_ _05055_ _05063_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ _04998_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10086_ _04915_ _04928_ _04953_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06388__I _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10131__C _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05903__A1 _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10988_ _00580_ clknet_leaf_13_clock exec.out_of_order_exec vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_206_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06459__A2 _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__I _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08908__A1 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08820_ _03207_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ _03860_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05963_ stack\[8\]\[4\] stack\[9\]\[4\] _01472_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10723__CLK clknet_leaf_50_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07702_ _02977_ _02972_ _02979_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05894_ _00820_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08682_ _03785_ _03809_ _03810_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ mem.mem_dff.code_mem\[30\]\[0\] _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05745__I1 stack\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07631__B _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07564_ _02869_ _02861_ _02872_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10873__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09097__B1 _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09303_ _04266_ _04286_ _04263_ _03624_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06515_ net242 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07647__A1 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07495_ _02816_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09234_ _04015_ _04109_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06446_ exec.memory_input\[7\] _01846_ _01976_ _01981_ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_167_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09165_ _04163_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_182_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06377_ _01816_ _01913_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08116_ _03308_ _03309_ _03310_ _03311_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07857__I _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input79_I rambus_wb_dat_i[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05328_ _00880_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09096_ _04119_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ _02985_ _02467_ _03248_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_123_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07078__B _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05259_ stack\[15\]\[0\] stack\[12\]\[0\] stack\[13\]\[0\] stack\[14\]\[0\] _00801_
+ _00803_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_163_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_21_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08375__A2 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09293__B _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06386__A1 stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10182__A2 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ _03007_ _04869_ _04876_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06386__B2 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08949_ _04015_ _04016_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06138__A1 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _00503_ clknet_leaf_141_clock stack\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10842_ _00434_ clknet_leaf_175_clock stack\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05361__A2 _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10237__A3 _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _00365_ clknet_leaf_53_clock net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08063__A1 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05287__I _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09982__I _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__B1 _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10746__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A2 _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10207_ _05046_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11187_ net243 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05424__I0 stack\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10138_ _04139_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05975__I1 stack\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10069_ _04932_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06129__A1 _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10896__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07007__I _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05951__S _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09079__B1 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__B1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06300_ _01191_ _01228_ _01237_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07280_ _02651_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06301__A1 _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06231_ _00838_ _01761_ _01236_ _01205_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_176_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06162_ _01113_ _01669_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06093_ _01636_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10400__A3 _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09921_ _04580_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06080__A3 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09003__B1 _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09852_ _04554_ _04767_ _04775_ net65 _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06368__A1 _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08803_ _03789_ _03901_ _03905_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09783_ _04413_ _01238_ _04725_ _04666_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06995_ mem.mem_dff.code_mem\[12\]\[4\] _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05966__I1 stack\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08109__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08734_ _03847_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05946_ _01278_ _01484_ _01487_ _01489_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05591__A2 stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07868__A1 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05877_ _01416_ _01418_ _01419_ _01420_ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08665_ _03235_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_215_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07616_ _02857_ _02905_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07361__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08596_ _03741_ _01685_ _01692_ _03640_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11051__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07547_ _02856_ _02848_ _02859_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09085__A3 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10619__CLK clknet_leaf_105_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07478_ mem.mem_dff.code_mem\[25\]\[5\] _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ _04208_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06429_ net151 _01716_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06491__I net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ stack\[1\]\[0\] _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output185_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10769__CLK clknet_leaf_31_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09079_ _04019_ _04110_ _04095_ _04112_ _04113_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05249__I3 stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11110_ _00702_ clknet_leaf_141_clock stack\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11041_ _00633_ clknet_leaf_34_clock cycles_per_ms\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06359__A1 _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07020__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05421__I3 stack\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _00417_ clknet_leaf_162_clock stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10756_ _00348_ clknet_leaf_48_clock mem.dff_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10091__A1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10687_ _00279_ clknet_leaf_61_clock mem.mem_dff.data_mem\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08036__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09784__A1 _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08587__A2 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09217__I _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05800_ _01258_ _01343_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06780_ _02255_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05731_ _01274_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11074__CLK clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__C _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _03620_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05662_ net258 _01197_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05480__I _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ mem.mem_dff.code_mem\[23\]\[4\] _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _03568_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05593_ _01062_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ _02688_ _02689_ _02691_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09887__I _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07263_ mem.mem_dff.code_mem\[19\]\[5\] _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10911__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09002_ _04045_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05884__I0 stack\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06214_ _01756_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07194_ _02557_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06017__S _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06145_ _01133_ _01671_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06076_ _01150_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09904_ _04596_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10137__A2 _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _04587_ _04762_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08031__I _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05939__I1 stack\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09766_ _04716_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05403__I3 stack\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ _02413_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08717_ _03217_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05929_ stack\[2\]\[3\] stack\[3\]\[3\] _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09697_ _04469_ _04470_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08502__A2 _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07091__B _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10441__CLK clknet_leaf_67_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08648_ _01763_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05390__I _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ _01891_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _00202_ clknet_leaf_92_clock mem.mem_dff.code_mem\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A1 mem.mem_dff.code_mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10591__CLK clknet_leaf_87_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _00133_ clknet_leaf_97_clock mem.mem_dff.code_mem\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05875__I0 stack\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08018__A1 _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _00064_ clknet_leaf_58_clock mem.mem_dff.code_mem\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08018__B2 stack\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08569__A2 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09465__C _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05565__I _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11024_ _00616_ clknet_leaf_17_clock cycles_per_ms\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__I _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05555__A2 stack\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05307__A2 _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__A2 _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10934__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_143_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ _00400_ clknet_leaf_163_clock stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10739_ _00331_ clknet_leaf_159_clock stack\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08009__A1 _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__B2 stack\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09757__A1 _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10367__A2 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput116 net116 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput127 net127 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput138 net138 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput149 net149 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10381__I stack\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07176__B _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ _02256_ _02989_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05794__A2 _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06901_ _02351_ _02352_ _02342_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_68_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07881_ _03090_ _03117_ _03113_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ delay_cycles\[5\] _04579_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06832_ _02264_ _02296_ _02283_ _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10464__CLK clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06743__A1 _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05546__A2 stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09551_ delay_cycles\[19\] _04510_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06763_ _02227_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _03238_ _03646_ _03657_ stack\[19\]\[6\] _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05714_ _00774_ _00766_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06694_ mem.mem_dff.code_mem\[4\]\[5\] _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09482_ _01697_ _04261_ _01668_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08433_ _03601_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05645_ _01188_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08364_ mem.mem_dff.code_mem\[5\]\[7\] _03352_ _03353_ mem.mem_dff.code_mem\[20\]\[7\]
+ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05576_ _01124_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _02677_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09996__A1 _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ mem.mem_dff.code_mem\[6\]\[5\] _03388_ _03389_ mem.mem_dff.code_mem\[30\]\[5\]
+ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ mem.mem_dff.code_mem\[19\]\[1\] _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__A1 _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ _02569_ _02564_ _02570_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10358__A2 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input61_I i_wb_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06128_ _01670_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08420__A1 _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08971__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06059_ _01599_ _01600_ _01602_ _01582_ _01064_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__05385__I _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09818_ _03737_ _04739_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08723__A2 _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06329__A4 _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__B _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09771__I1 _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ _03619_ _04277_ _04705_ _04467_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10957__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 i_wb_addr[0] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_122_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05848__I0 stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10524_ _00116_ clknet_leaf_110_clock mem.mem_dff.code_mem\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput29 i_wb_addr[1] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09739__A1 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _00047_ clknet_leaf_70_clock mem.mem_dff.code_mem\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10386_ _03218_ _05172_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08175__C2 _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11007_ _00599_ clknet_leaf_13_clock prev_level_interrupt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09762__I1 _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06120__S _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07015__I _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10285__A1 _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05430_ _00981_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06854__I _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__CLK clknet_leaf_178_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05361_ _00889_ _00911_ _00913_ _00878_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10376__I _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _02508_ _02501_ _02509_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08080_ net117 _03272_ _03278_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05292_ _00789_ _00845_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08650__A1 _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07031_ mem.mem_dff.code_mem\[13\]\[4\] _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09386__B _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08402__A1 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05216__A1 _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08953__A2 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05419__B _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08982_ _04038_ _04039_ _04041_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05767__A2 stack\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__S1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ mem.mem_dff.data_mem\[6\]\[2\] _03156_ _03152_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07864_ _02036_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09603_ _04545_ _04533_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06815_ _02282_ _02274_ _02283_ _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07795_ _03051_ _03046_ _03052_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06192__A2 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ delay_cycles\[17\] delay_cycles\[16\] _04493_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06746_ _02227_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__A1 _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09130__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09465_ _04371_ _04433_ _04434_ _04324_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06677_ _02102_ _02176_ _02166_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08416_ net126 _03122_ _03591_ _03592_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_40_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05628_ _01173_ _01174_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09396_ _04369_ _04370_ _04372_ _04266_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10028__B2 _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08347_ mem.mem_dff.data_mem\[0\]\[6\] _03475_ _03476_ _03536_ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05559_ _01083_ stack\[24\]\[6\] stack\[25\]\[6\] _01078_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08278_ mem.mem_dff.code_mem\[9\]\[4\] _03429_ _03430_ mem.mem_dff.code_mem\[28\]\[4\]
+ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05455__A1 _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05455__B2 stack\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07229_ _02523_ _02605_ _02600_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07595__I mem.mem_dff.code_mem\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__A2 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _01715_ _03990_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ _04998_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06955__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06939__I _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06707__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06183__A2 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09050__I _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10019__A1 delay_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05694__A1 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09985__I _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08632__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _00099_ clknet_leaf_111_clock mem.mem_dff.code_mem\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07986__A3 _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05997__A2 _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _00030_ clknet_leaf_75_clock mem.mem_dff.code_mem\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06115__S net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07199__A1 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08935__A2 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _05066_ _05165_ _05166_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08699__A1 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07371__A1 _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06174__A2 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06600_ _02045_ _02103_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ mem.mem_dff.code_mem\[28\]\[3\] _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10258__A1 _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _02054_ _02049_ _02057_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10258__B2 _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10502__CLK clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06584__I _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09250_ _04220_ _04236_ _04238_ stack\[22\]\[2\] _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_209_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _01622_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08871__A1 _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08871__B2 stack\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08201_ mem.mem_dff.code_mem\[8\]\[2\] _02293_ _02701_ mem.mem_dff.code_mem\[22\]\[2\]
+ _03394_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05413_ _00963_ _00927_ stack\[22\]\[3\] _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09181_ stack\[20\]\[0\] _04189_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06393_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__CLK clknet_leaf_94_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08132_ _03098_ _03042_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05344_ _00889_ _00893_ _00896_ _00878_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_147_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05437__A1 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05437__B2 _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08063_ net114 _03250_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05275_ _00825_ _00826_ _00829_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _02441_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09179__A2 _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11008__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08926__A2 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08965_ _04024_ _04028_ _04030_ stack\[0\]\[0\] _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ mem.mem_dff.data_mem\[5\]\[5\] _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08896_ _03819_ _03970_ _03977_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input24_I i_wb_addr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _02978_ _03087_ _03082_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ _03010_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _04249_ _01623_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09103__A2 _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06729_ mem.mem_dff.code_mem\[5\]\[5\] _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ _01891_ _04380_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08862__A1 _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _04298_ _04356_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08614__A1 stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05428__B2 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06443__B _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10223_ _04225_ _05045_ _05062_ stack\[12\]\[4\] _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06928__A1 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05774__S _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10154_ _05007_ _05009_ _05010_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_216_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05600__A1 _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10085_ _04940_ _04942_ _04947_ _04952_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05573__I _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09045__I _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A1 _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07105__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10987_ _00579_ clknet_leaf_39_clock mem.mem_io.past_write vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08302__B1 _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10675__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05419__A1 _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06092__A1 _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__B1 _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08369__C2 _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08908__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09030__A1 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07963__I _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05278__S0 _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _03859_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05962_ stack\[10\]\[4\] stack\[11\]\[4\] _01417_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05483__I _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_173_clock clknet_4_1_0_clock clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07701_ _02978_ _02973_ _02969_ _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08681_ _03650_ _03805_ _03803_ stack\[5\]\[1\] _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07344__A1 _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _01408_ _01431_ _01435_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07632_ _02922_ _02915_ _02924_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07563_ _02870_ _02862_ _02871_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_188_clock clknet_4_1_0_clock clknet_leaf_188_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09097__B2 stack\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ mem.io_data_out\[1\] _04285_ _03242_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06514_ mem.mem_dff.code_mem\[0\]\[3\] _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07494_ _02030_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A1 _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_191_clock_I clknet_4_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _04180_ _04208_ _04228_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ _01226_ _01977_ _01978_ _01980_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xclkbuf_leaf_111_clock clknet_4_13_0_clock clknet_leaf_111_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ _03721_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06376_ _01122_ _01745_ _01779_ _01026_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08115_ mem.mem_dff.code_mem\[3\]\[0\] _02136_ _02172_ mem.mem_dff.code_mem\[4\]\[0\]
+ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05327_ _00785_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09095_ _01856_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06083__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _03249_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05258_ _00789_ _00812_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05269__S0 _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10548__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09997_ _04870_ _01949_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06386__A2 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _03230_ _03848_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05393__I _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output130_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output228_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _01963_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_218_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__B1 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ _00502_ clknet_leaf_179_clock stack\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10698__CLK clknet_leaf_62_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07886__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _00433_ clknet_leaf_176_clock stack\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09088__A1 _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10772_ _00364_ clknet_leaf_53_clock net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A1 stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__A4 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05649__A1 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06310__A2 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09260__A1 stack\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__B2 stack\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08879__I _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06901__B _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10206_ _05045_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_90_clock clknet_4_15_0_clock clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08220__C1 mem.mem_dff.data_mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11186_ net245 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05424__I1 stack\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _04993_ _04995_ _04997_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06399__I _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10068_ net34 _04922_ _04929_ _04930_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__07326__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07732__B _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__B2 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06301__A2 _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06230_ _01205_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_clock clknet_4_3_0_clock clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06161_ _01699_ _01703_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_157_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__A1 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05478__I _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A1 _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06092_ _01633_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05812__A1 _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09003__A1 _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05812__B2 _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__B2 stack\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07693__I _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_clock clknet_4_14_0_clock clknet_leaf_58_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09851_ _04374_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_138_clock_I clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06368__A2 _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _03839_ _03899_ _03903_ stack\[6\]\[3\] _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _01224_ _01245_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06994_ _02424_ _02417_ _02426_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10840__CLK clknet_leaf_177_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _01931_ _03848_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05945_ _01485_ stack\[22\]\[4\] _01298_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_39_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08664_ _01926_ _03230_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05876_ _01271_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05718__I2 stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05941__I _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09413__I _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07615_ _02897_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08457__C _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05879__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08595_ _01676_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10990__CLK clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ _02857_ _02849_ _02858_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08029__I _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08817__A1 _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07477_ _02801_ _02802_ _02804_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input91_I rambus_wb_dat_i[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _01182_ _04208_ _04214_ _04216_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06428_ stack\[2\]\[6\] _01718_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05500__B1 _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10294__I _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _04163_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08045__A2 _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06359_ _01865_ _01871_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05388__I _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06056__A1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09078_ stack\[23\]\[7\] _04096_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output178_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _03234_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _00632_ clknet_leaf_34_clock cycles_per_ms\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08753__B1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07108__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07308__A1 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10824_ _00416_ clknet_leaf_162_clock stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10755_ _00347_ clknet_leaf_48_clock mem.dff_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10686_ _00278_ clknet_leaf_62_clock mem.mem_dff.data_mem\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09233__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07727__B _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05962__S _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05730_ _00805_ _01270_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_209_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__C _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05661_ _01188_ _01198_ _01200_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07400_ _02741_ _02733_ _02744_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08380_ _02003_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05592_ _01094_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07331_ _02604_ _02690_ _02686_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08275__A2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_64_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06286__A1 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07262_ _02634_ _02635_ _02637_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05333__I0 stack\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09001_ _03716_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06213_ _01720_ _01727_ _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05884__I1 stack\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07193_ mem.mem_dff.code_mem\[17\]\[7\] _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06144_ _01127_ _01670_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06589__A2 _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08983__B1 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06075_ _01583_ _01591_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _04810_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07538__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09834_ _04299_ _04758_ _04764_ _04761_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09765_ exec.memory_input\[2\] _04297_ _04715_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06977_ _02287_ _02412_ _02171_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08716_ _03785_ _03826_ _03836_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06767__I _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05928_ _00899_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _04640_ _04645_ _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08187__C _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08647_ _01183_ _03775_ _03784_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05859_ _00809_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08578_ _03707_ _03726_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07529_ _02022_ _02318_ _02133_ _02618_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_168_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10540_ _00132_ clknet_leaf_98_clock mem.mem_dff.code_mem\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05875__I1 stack\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _00063_ clknet_leaf_58_clock mem.mem_dff.code_mem\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09215__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08018__A2 _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06029__A1 _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__B1 _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09318__I _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05846__I _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11023_ _00615_ clknet_leaf_16_clock cycles_per_ms\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07282__B _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05581__I _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__B1 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__I0 stack\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10807_ _00399_ clknet_leaf_140_clock stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09454__A1 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10738_ _00330_ clknet_leaf_65_clock mem.mem_dff.data_mem\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09206__A1 _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08009__A2 _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10669_ _00261_ clknet_leaf_59_clock mem.mem_dff.code_mem\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput117 net117 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08965__B1 _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput128 net128 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput139 net139 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_177_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__I _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06440__A1 _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06440__B2 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__CLK clknet_leaf_34_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06900_ _02348_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ mem.mem_dff.data_mem\[4\]\[5\] _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10609__CLK clknet_leaf_92_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08193__B2 mem.mem_dff.code_mem\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ mem.mem_dff.code_mem\[8\]\[1\] _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06743__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09550_ delay_cycles\[18\] delay_cycles\[17\] _04509_ _04493_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06587__I _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06762_ _02116_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05491__I _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__B1 _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08501_ _03662_ _03664_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05713_ _00778_ _01256_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10759__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ _04439_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06693_ _02185_ _02186_ _02188_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09693__A1 _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__A2 _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08432_ _02045_ _03602_ _03608_ _03605_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07920__B _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05644_ _01184_ _01186_ _01187_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ mem.mem_dff.code_mem\[1\]\[7\] _02071_ _02562_ mem.mem_dff.code_mem\[17\]\[7\]
+ _02027_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08248__A2 _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05575_ _01123_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07314_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10055__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ mem.mem_dff.code_mem\[15\]\[5\] _03368_ _03369_ mem.mem_dff.code_mem\[29\]\[5\]
+ _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09996__A2 _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07211__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07245_ _02617_ _02622_ _02624_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05867__S _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09748__A2 _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ _02478_ _02565_ _02558_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07367__B _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06271__B _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I i_wb_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06431__A1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _01581_ _01601_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09817_ net190 _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06497__I _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05793__I0 stack\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09748_ _03625_ _01241_ intr\[0\] _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output210_I net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _04500_ _04501_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09684__A1 _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07830__B _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07121__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10523_ _00115_ clknet_leaf_110_clock mem.mem_dff.code_mem\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 i_wb_addr[10] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05848__I1 stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10454_ _00046_ clknet_leaf_71_clock mem.mem_dff.code_mem\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09739__A2 _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10385_ stack\[15\]\[2\] _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05576__I _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05225__A2 _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_12_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08175__B2 mem.mem_dff.code_mem\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ _00598_ clknet_leaf_12_clock single_step vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10901__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06200__I _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06489__A1 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10285__A2 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08127__I _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09978__A2 _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05360_ _00894_ _00905_ _00912_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07989__A1 _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05291_ stack\[19\]\[1\] stack\[16\]\[1\] stack\[17\]\[1\] stack\[18\]\[1\] _00843_
+ _00844_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08650__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07030_ _02452_ _02445_ _02454_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08402__A2 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10431__CLK clknet_leaf_76_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05486__I _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05216__A2 _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A1 _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08981_ _04040_ _04021_ _04035_ stack\[0\]\[6\] _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07932_ _02994_ _03155_ _03158_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06016__I1 stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ mem.mem_dff.data_mem\[4\]\[1\] _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06814_ _02251_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09602_ _04559_ _04561_ _04558_ cycles_per_ms\[8\] _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07794_ _02936_ _03047_ _03039_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09533_ _04486_ _04487_ _04488_ _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_06745_ _02101_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08469__A2 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09464_ _03737_ _04380_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05790__I3 stack\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06676_ _02174_ _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09421__I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08415_ net126 _03588_ _03589_ _03122_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ net190 net189 _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09395_ _03889_ _04371_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09418__A1 _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08346_ _03533_ _03534_ _03535_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10028__A2 _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05558_ _01103_ _01104_ _01106_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ mem.mem_dff.code_mem\[16\]\[4\] _02536_ _03463_ _03468_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05489_ _01028_ _01032_ _01035_ _01038_ _00920_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_153_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06652__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ mem.mem_dff.code_mem\[18\]\[6\] _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05455__A2 stack\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ mem.mem_dff.code_mem\[16\]\[7\] _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06404__A1 _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output160_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10170_ _05019_ _05021_ _05022_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06955__A2 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10924__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_186_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__I _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06707__A2 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07116__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09409__A1 _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06904__B _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06690__I _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10506_ _00098_ clknet_leaf_109_clock mem.mem_dff.code_mem\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _00029_ clknet_leaf_73_clock mem.mem_dff.code_mem\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07199__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08396__A1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10368_ _05068_ _05155_ _05161_ stack\[17\]\[6\] _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07735__B _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ _05111_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__A1 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05757__I0 stack\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06174__A3 _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09648__A1 _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _02056_ _02052_ _02046_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10258__A2 _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05509__I0 stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09241__I _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08320__A1 _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06461_ mem.mem_dff.cycles\[1\] mem.mem_dff.cycles\[0\] _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08871__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _03387_ _03390_ _03393_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05412_ _00927_ stack\[20\]\[3\] stack\[21\]\[3\] _00963_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09180_ _04188_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05685__A2 _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06392_ _01928_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08131_ _03043_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05343_ _00894_ _00826_ _00895_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__I mem.mem_dff.code_mem\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05437__A2 stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ net71 _03252_ _03254_ net122 _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05274_ stack\[27\]\[0\] stack\[24\]\[0\] stack\[25\]\[0\] stack\[26\]\[0\] _00827_
+ _00828_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07013_ _02345_ _02440_ _02198_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_175_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09844__C _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08964_ _04029_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08139__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09336__B1 _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _03143_ _03144_ _03146_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08895_ _03776_ _03972_ _03976_ stack\[10\]\[0\] _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_151_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07846_ mem.mem_dff.data_mem\[3\]\[6\] _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I i_la_write vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07777_ mem.mem_dff.data_mem\[1\]\[7\] _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06728_ _02212_ _02213_ _02215_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06775__I _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09516_ _04249_ _04251_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08311__A1 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09447_ _04417_ _04405_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06659_ _02160_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05612__C _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08862__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10477__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08990__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05676__A2 _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09378_ _04354_ net64 _04355_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05920__I0 stack\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08329_ _03518_ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08075__B1 _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09811__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08614__A2 _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05279__I2 stack\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10222_ _05047_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07050__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10153_ _04288_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11102__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05854__I _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10084_ _04629_ _04950_ _04951_ intr_enable\[0\] _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A1 _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__B2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05739__I0 stack\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06156__A3 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10986_ _00578_ clknet_leaf_9_clock net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05911__I0 stack\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08605__A2 _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__I _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06092__A2 _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08369__B2 mem.mem_dff.code_mem\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__S _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__A1 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09030__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05278__S1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05978__I0 stack\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08140__I _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I i_la_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05961_ _01480_ _01500_ _01502_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_140_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09869__A1 _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ _02059_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09869__B2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08680_ _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05892_ _01305_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07344__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07631_ _02870_ _02916_ _02923_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06595__I _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07562_ _02841_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09097__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ _04282_ _04284_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06513_ _02039_ _02029_ _02042_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _02816_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10100__A1 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_134_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _04227_ _04210_ _04223_ stack\[21\]\[5\] _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06855__A1 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06444_ _01968_ _01979_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09163_ _04175_ _04171_ _04176_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06375_ exec.memory_input\[5\] _01744_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08114_ mem.mem_dff.code_mem\[19\]\[0\] _02619_ _02675_ mem.mem_dff.code_mem\[21\]\[0\]
+ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06607__A1 _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05326_ _00878_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09094_ _04054_ _04115_ _04125_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _02985_ _02256_ _03248_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__06083__A2 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05257_ stack\[11\]\[0\] stack\[8\]\[0\] stack\[9\]\[0\] stack\[10\]\[0\] _00811_
+ _00794_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11125__CLK clknet_leaf_158_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05875__S _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05269__S1 _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09996_ _04866_ _01904_ _04875_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05674__I _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07583__A2 _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_59_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__I _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05594__A1 stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ _03691_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05594__B2 stack\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _03961_ _03942_ _03962_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__B2 stack\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output123_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07829_ _02040_ _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10840_ _00432_ clknet_leaf_177_clock stack\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09088__A2 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07099__A1 _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _00363_ clknet_leaf_53_clock net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__A2 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05649__A2 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__C _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09260__A2 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10158__A1 _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__A2 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ stack\[12\]\[0\] _05048_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07285__B _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11185_ net247 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08771__A1 _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ net182 _04996_ _03183_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05424__I2 stack\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10067_ _04934_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10642__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__A1 _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08523__B2 stack\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _00561_ clknet_4_3_0_clock net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11148__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ _01701_ _01702_ _01648_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10397__A1 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A2 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _01634_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07974__I _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A2 _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ _04774_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A1 _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08801_ _03787_ _03901_ _03904_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_60_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06993_ _02394_ _02418_ _02425_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09781_ _04723_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05944_ _00900_ stack\[23\]\[4\] _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08732_ _03636_ _01925_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A1 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08663_ _03794_ _03774_ _03795_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05875_ stack\[30\]\[6\] stack\[31\]\[6\] _01360_ _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10321__A1 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05718__I3 stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07614_ mem.mem_dff.code_mem\[29\]\[3\] _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05879__A2 _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08594_ _02002_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07214__I mem.mem_dff.code_mem\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07545_ _02841_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08817__A2 _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_12_0_clock clknet_3_6_0_clock clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07476_ _02717_ _02803_ _02799_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A2 _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09215_ _03898_ _04215_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06427_ _01963_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05500__A1 stack\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05500__B2 stack\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _04071_ _04161_ _04162_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input84_I rambus_wb_dat_i[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06358_ _01722_ net62 _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_202_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10515__CLK clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05309_ stack\[3\]\[1\] stack\[0\]\[1\] stack\[1\]\[1\] stack\[2\]\[1\] _00811_ _00794_
+ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_198_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _03855_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06289_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07884__I _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _03233_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08753__A1 _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08753__B2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05567__A1 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _03627_ _04864_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08505__A1 _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09702__B1 _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10312__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08269__B1 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10823_ _00415_ clknet_leaf_160_clock stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06119__I0 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10754_ _00346_ clknet_leaf_42_clock mem.io_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _00277_ clknet_leaf_60_clock mem.mem_dff.data_mem\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05342__I1 stack\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05579__I _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09233__A2 _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10379__A1 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07244__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06047__A2 _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05350__S0 _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_187_clock clknet_4_1_0_clock clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08339__A4 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_110_clock clknet_4_13_0_clock clknet_leaf_110_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10119_ _04956_ _04981_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__B _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11099_ _00691_ clknet_leaf_32_clock net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10303__A1 stack\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05660_ _01195_ _01203_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_125_clock clknet_4_12_0_clock clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05591_ _01130_ stack\[12\]\[7\] stack\[13\]\[7\] _01131_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05730__A1 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ _02677_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10538__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _02604_ _02636_ _02632_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06286__A2 _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05333__I1 stack\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ _04054_ _04052_ _04055_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05494__B1 stack\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06212_ _01197_ _01737_ _01753_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07192_ _02580_ _02575_ _02581_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ _01597_ _01621_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10688__CLK clknet_leaf_61_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__B2 stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06074_ _01617_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _04805_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09833_ _04603_ _04762_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05549__A1 _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09852__C _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09764_ _04711_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06976_ _02318_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ _03835_ _03830_ _03833_ stack\[8\]\[1\] _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05927_ _01380_ _01466_ _01470_ _01436_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09695_ _04646_ _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__A1 _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ stack\[20\]\[6\] stack\[21\]\[6\] _00810_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08646_ _03776_ _03779_ _03783_ stack\[4\]\[0\] _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05789_ _01282_ _01325_ _01332_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08577_ _01999_ _03699_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ mem.mem_dff.code_mem\[27\]\[0\] _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07459_ _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output190_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10470_ _00062_ clknet_leaf_57_clock mem.mem_dff.code_mem\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09215__A2 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05580__S0 _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07226__A1 _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _04124_ _04147_ _04149_ stack\[18\]\[2\] _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__B2 stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05332__S0 _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ _00614_ clknet_leaf_15_clock cycles_per_ms\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08726__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07563__B _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05960__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_clock clknet_4_9_0_clock clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__B2 _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05399__S0 _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05712__A1 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05563__I1 stack\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10806_ _00398_ clknet_leaf_134_clock stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_57_clock clknet_4_14_0_clock clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06268__A2 _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _00329_ clknet_leaf_65_clock mem.mem_dff.data_mem\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08662__B1 _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10830__CLK clknet_leaf_153_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _00260_ clknet_leaf_55_clock mem.mem_dff.code_mem\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09206__A2 _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07738__B _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_2_0_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10599_ _00191_ clknet_leaf_100_clock mem.mem_dff.code_mem\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09509__I _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A1 _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08965__B2 stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput118 net118 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput129 net129 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09765__I0 exec.memory_input\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06830_ _02285_ _02295_ _02297_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06761_ _02227_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08500_ _03663_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05712_ _01255_ _01087_ _01105_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09142__B2 stack\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06692_ _02117_ _02187_ _02183_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09480_ _01131_ _04439_ _04447_ _04448_ _04401_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09693__A2 _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ net115 _03603_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05643_ net134 net133 _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05703__A1 _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__I mem.mem_dff.code_mem\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08362_ mem.mem_dff.code_mem\[16\]\[7\] _02536_ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05574_ _01122_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07313_ _02648_ _02676_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06259__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08293_ _03484_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10055__A3 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07244_ _02591_ _02623_ _02615_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07208__A1 _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07175_ mem.mem_dff.code_mem\[17\]\[2\] _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _00699_ _01668_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06057_ _01114_ _01583_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input47_I i_wb_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09816_ _04749_ _04744_ _04750_ _04751_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09747_ _04685_ _04659_ _04704_ _02010_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ _02384_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05942__A1 _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05615__C _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05793__I1 stack\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10279__B1 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08993__I _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _04505_ _04504_ _04624_ _04636_ _04637_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ _03732_ _03767_ _03768_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output203_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06727__B _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10853__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__I _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_182_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__A1 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11071__D _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10522_ _00114_ clknet_leaf_112_clock mem.mem_dff.code_mem\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09757__C _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ _00045_ clknet_leaf_73_clock mem.mem_dff.code_mem\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09739__A3 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05857__I _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10384_ _05176_ _05171_ _05177_ _05178_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05305__S0 _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06422__A2 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05793__S _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11005_ _00597_ clknet_leaf_128_clock exec.memory_input\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06186__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05592__I _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09064__I _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09675__A2 _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06489__A2 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05541__B _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08408__I _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07312__I _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10159__B _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A2 _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05290_ _00793_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06413__A2 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _03237_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__I _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07931_ mem.mem_dff.data_mem\[6\]\[1\] _03156_ _03152_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10726__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08166__A2 _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A1 _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06598__I mem.mem_dff.code_mem\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03097_ _03103_ _03105_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ delay_cycles\[9\] _04560_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06813_ _02164_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07793_ mem.mem_dff.data_mem\[2\]\[2\] _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09532_ delay_cycles\[12\] delay_cycles\[11\] delay_cycles\[10\] _04491_ _04492_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06744_ _02227_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07931__B _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10876__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06675_ _02174_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07677__A1 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _04431_ _04432_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08874__B1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input101_I rambus_wb_dat_i[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ _03594_ _03595_ _03596_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05626_ net188 _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09394_ _04367_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07429__A1 _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08345_ mem.mem_dff.data_mem\[4\]\[6\] _03323_ _03324_ mem.mem_dff.data_mem\[5\]\[6\]
+ _03325_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05557_ stack\[30\]\[6\] _01105_ _01076_ stack\[31\]\[6\] _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08276_ _03464_ _03465_ _03466_ _03467_ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05488_ _01028_ _01037_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06101__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07227_ _02607_ _02603_ _02609_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08929__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09149__I _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07158_ _02554_ _02549_ _02555_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06109_ net110 _01629_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07089_ _02500_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output153_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05345__C _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09106__A1 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09657__A2 _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09121__A4 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09409__A2 _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A1 _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11031__CLK clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08093__A1 _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _00097_ clknet_leaf_106_clock mem.mem_dff.code_mem\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07288__B _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__A1 _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _00028_ clknet_leaf_74_clock mem.mem_dff.code_mem\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09042__B1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10749__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08396__A2 _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10367_ _03662_ _03692_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05603__B1 stack\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _03870_ _03941_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09345__A1 _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06159__A1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10899__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07307__I _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05906__A1 _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05757__I1 stack\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A2 _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10112__C1 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06367__B _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06460_ _01994_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07042__I mem.mem_dff.code_mem\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05411_ _00962_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08608__B1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06391_ _01679_ _01686_ _01927_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08130_ mem.mem_dff.data_mem\[4\]\[0\] _03323_ _03324_ mem.mem_dff.data_mem\[5\]\[0\]
+ _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07977__I _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05342_ stack\[23\]\[2\] stack\[20\]\[2\] stack\[21\]\[2\] stack\[22\]\[2\] _00822_
+ _00823_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05517__S0 _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09820__A2 _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08061_ _03262_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05273_ _00784_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07012_ _02318_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05842__B1 _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06398__A1 _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ _03973_ _04027_ _04021_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09336__A1 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07914_ _03086_ _03145_ _03141_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09336__B2 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ _03975_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07845_ _03089_ _03085_ _03091_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07661__B _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07776_ _03036_ _03031_ _03037_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11054__CLK clknet_leaf_25_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ _04299_ _04475_ _04476_ _04467_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06727_ _02117_ _02214_ _02210_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08847__B1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08048__I _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06658_ net235 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_209_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05609_ _01137_ _01156_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_185_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09377_ _04354_ _01986_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06589_ _02094_ _02100_ _02104_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__B1 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08075__A1 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08328_ mem.mem_dff.code_mem\[10\]\[6\] _03343_ _03344_ mem.mem_dff.code_mem\[24\]\[6\]
+ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08075__B2 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08259_ _03289_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05279__I3 stack\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05833__B1 _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09575__A1 delay_cycles\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10221_ _03721_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _04610_ _05008_ _05001_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08511__I _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09327__A1 _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _04936_ _04945_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07127__I _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06031__I _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06966__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06561__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05870__I _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09342__I _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _00577_ clknet_leaf_131_clock net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10421__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06313__A1 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10571__CLK clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09015__B1 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08369__A2 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _00011_ clknet_leaf_122_clock mem.mem_dff.code_mem\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__A2 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07041__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05978__I1 stack\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05960_ _01398_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09869__A2 _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05981__S _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05891_ _01416_ _01432_ _01433_ _01434_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07630_ _02897_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07561_ _02526_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08829__B1 _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09300_ _04283_ mem.dff_data_out\[1\] _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06512_ _02041_ _02032_ _02033_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _02759_ _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06304__A1 _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10100__A2 _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ _01922_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06855__A2 _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06443_ _01975_ _01732_ _01635_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08057__A1 mem.io_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09162_ _04126_ _04166_ _04164_ stack\[1\]\[3\] _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06374_ _01898_ _01911_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ mem.mem_dff.code_mem\[2\]\[0\] _02097_ _02587_ mem.mem_dff.code_mem\[18\]\[0\]
+ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05325_ _00806_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09093_ _04124_ _04117_ _04120_ stack\[24\]\[2\] _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08044_ _03247_ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09006__B1 _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05256_ _00810_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05418__I0 stack\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09427__I _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09995_ _02056_ _04867_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _03961_ _03992_ _04014_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _03844_ _03946_ _03955_ stack\[26\]\[5\] _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_218_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08532__A2 _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07828_ mem.mem_dff.data_mem\[3\]\[2\] _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07759_ mem.mem_dff.data_mem\[1\]\[2\] _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output116_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08296__A1 mem.mem_dff.code_mem\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _00362_ clknet_leaf_31_clock net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__B2 mem.mem_dff.code_mem\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10594__CLK clknet_leaf_90_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _03621_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__A2 _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10204_ _05047_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07023__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08220__B2 mem.mem_dff.data_mem\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11184_ net250 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10135_ _04955_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08771__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10066_ net34 _04929_ _04930_ _04933_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_48_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09720__A1 _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05533__C _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10968_ _00560_ clknet_leaf_43_clock net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09800__I _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10899_ _00491_ clknet_leaf_186_clock stack\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ _01251_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _03837_ _03899_ _03903_ stack\[6\]\[2\] _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__A2 _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10467__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _04412_ _04477_ _03620_ _02127_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ _02377_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07990__I _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _03234_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05943_ _01485_ stack\[20\]\[4\] _01303_ _01486_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09711__A1 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05724__B _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ _03659_ _03778_ _03792_ stack\[4\]\[5\] _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06525__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05874_ stack\[28\]\[6\] stack\[29\]\[6\] _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05959__S0 _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10321__A2 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _02909_ _02904_ _02910_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08593_ _03736_ _03704_ _03739_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07544_ _02511_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07475_ _02790_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09214_ _04210_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06426_ _01962_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05500__A2 _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09778__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09145_ _01617_ _03679_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06357_ _01767_ _01894_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09242__A3 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10388__A2 _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input77_I rambus_wb_ack_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05308_ _00846_ _00849_ _00854_ _00861_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09076_ _04038_ _04110_ _04111_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06288_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _03190_ _01711_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05239_ _00793_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08061__I _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08753__A2 _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09978_ delay_cycles\[23\] _04810_ _04859_ _04499_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06764__A1 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08929_ _03890_ _03992_ _04000_ _04002_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09702__A1 _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05634__B _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09702__B2 _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10312__A2 _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ _00414_ clknet_leaf_161_clock stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06119__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ _00345_ clknet_leaf_41_clock mem.io_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _00276_ clknet_leaf_62_clock mem.mem_dff.data_mem\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07492__A2 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05342__I2 stack\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10379__A2 _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05796__S _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08441__A1 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06047__A3 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08292__I1 _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09495__C _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05350__S1 _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__A1 _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__I _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_177_clock_I clknet_4_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05802__I0 stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _04593_ _04963_ _04944_ _00778_ _04406_ _04939_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11098_ _00690_ clknet_leaf_14_clock net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ net22 net21 net24 net23 _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__06507__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10303__A2 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07180__A1 _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11115__CLK clknet_leaf_192_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05590_ _01127_ _01128_ _01136_ _01137_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05730__A2 _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__I0 stack\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _02621_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08146__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05333__I2 stack\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05494__A1 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06211_ _01719_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07191_ _02523_ _02576_ _02572_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05494__B2 _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01684_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08432__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08983__A2 _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06073_ _01588_ _01605_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_172_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ _04598_ _04806_ _04809_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08196__B1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _03623_ _04758_ _04763_ _04761_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09763_ _04714_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06975_ _02017_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08714_ _03214_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05926_ _01467_ _01468_ _01469_ _01434_ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09694_ _04254_ _04477_ _04649_ _04652_ _04653_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07225__I _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09160__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05857_ _01266_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08257__S _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08576_ _03724_ _03711_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05721__A2 _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05788_ _01299_ _01328_ _01331_ _01304_ _01275_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07527_ _02839_ _02830_ _02843_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07458_ _02759_ _02789_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05485__A1 _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ _01905_ _01944_ _01941_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ mem.mem_dff.code_mem\[23\]\[1\] _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07895__I _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05580__S1 _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10632__CLK clknet_leaf_115_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _04050_ _04144_ _04151_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output183_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09059_ stack\[23\]\[2\] _04090_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08974__A2 _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05332__S1 _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11069__D _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10782__CLK clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _00613_ clknet_leaf_16_clock cycles_per_ms\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08726__A2 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__B _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06737__A1 _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11138__CLK clknet_leaf_187_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09151__A2 _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07162__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05399__S1 _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05712__A2 _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10049__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05563__I2 stack\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _00397_ clknet_leaf_139_clock stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10736_ _00328_ clknet_leaf_65_clock mem.mem_dff.data_mem\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08662__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10667_ _00259_ clknet_leaf_55_clock mem.mem_dff.code_mem\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07217__A2 _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08414__A1 _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10598_ _00190_ clknet_leaf_99_clock mem.mem_dff.code_mem\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08965__A2 _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput119 net119 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__I _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_6_0_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__I1 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07754__B _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06760_ mem.mem_dff.code_mem\[6\]\[4\] _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09142__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__A1 _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05711_ _00773_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10505__CLK clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06691_ _02174_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08430_ _02041_ _03602_ _03607_ _03605_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05642_ _01185_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08361_ _03544_ _03547_ _03548_ _03549_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05573_ _01121_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08102__B1 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07312_ _02675_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10655__CLK clknet_leaf_95_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07456__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ mem.dff_data_out\[4\] _03482_ _03483_ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__A1 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10055__A4 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05467__A1 stack\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _02621_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05467__B2 stack\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07929__B _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ _02567_ _02564_ _02568_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ prev_reg_write _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_219_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06967__A1 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ _01574_ _01232_ _01064_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09863__C _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07664__B _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _04423_ _04730_ _04724_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10090__B _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09746_ _04403_ _04656_ _04703_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06958_ _02384_ _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_171_clock clknet_4_3_0_clock clknet_leaf_171_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05942__A2 stack\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09133__A2 _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10279__A1 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05909_ _01401_ _01451_ _01452_ _01405_ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10279__B2 stack\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _04625_ _04626_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _02314_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _03694_ _03763_ _03760_ stack\[3\]\[6\] _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08892__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_186_clock clknet_4_1_0_clock clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08559_ _03707_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_125_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _00113_ clknet_leaf_112_clock mem.mem_dff.code_mem\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10452_ _00044_ clknet_leaf_72_clock mem.mem_dff.code_mem\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09739__A4 _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10383_ net145 _05174_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05305__S1 _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06034__I _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_124_clock clknet_4_12_0_clock clknet_leaf_124_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05630__A1 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11004_ _00596_ clknet_leaf_129_clock exec.memory_input\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10528__CLK clknet_leaf_113_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05806__C _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_139_clock clknet_4_7_0_clock clknet_leaf_139_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08332__B1 _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10678__CLK clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A1 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A1 _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05449__A1 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10719_ _00311_ clknet_leaf_30_clock mem.mem_dff.data_mem\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10175__B _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ _02984_ _03155_ _03157_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06879__I _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09363__A2 mem.dff_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ _03073_ _03104_ _03095_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07374__A1 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09600_ _04555_ _04556_ _04490_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06812_ mem.mem_dff.code_mem\[7\]\[7\] _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07792_ _03049_ _03046_ _03050_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ delay_cycles\[9\] delay_cycles\[8\] delay_cycles\[7\] _04490_ _04491_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06743_ _02169_ _02226_ _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09462_ net156 net155 _04405_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_92_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06674_ _02169_ _02173_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08874__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10130__B1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08874__B2 stack\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08413_ net125 _02121_ _03591_ _03592_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05625_ mem.sram_enable _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09393_ exec.out_of_order_exec _04359_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_178_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08344_ mem.mem_dff.data_mem\[1\]\[6\] _03015_ _03069_ mem.mem_dff.data_mem\[3\]\[6\]
+ mem.mem_dff.data_mem\[7\]\[6\] _03379_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_05556_ _01045_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08275_ mem.mem_dff.code_mem\[3\]\[4\] _03364_ _03365_ mem.mem_dff.code_mem\[4\]\[4\]
+ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05487_ _01036_ stack\[19\]\[5\] _01033_ stack\[18\]\[5\] _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06101__A2 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ _02608_ _02605_ _02600_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_41_clock clknet_4_9_0_clock clknet_leaf_41_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08929__A2 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ _02523_ _02550_ _02546_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06108_ _01633_ _01646_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07601__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _02411_ _02499_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06039_ _01252_ _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06789__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_56_clock clknet_4_12_0_clock clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_51_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__A2 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10820__CLK clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09106__A2 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04667_ _04687_ _04673_ _04324_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08314__B1 _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__S _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08509__I _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08865__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07413__I mem.mem_dff.code_mem\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10970__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A2 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__A1 mem.io_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ _00096_ clknet_leaf_109_clock mem.mem_dff.code_mem\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05851__A1 _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _00027_ clknet_leaf_73_clock mem.mem_dff.code_mem\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05851__B2 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09042__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09042__B2 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_7_0_clock clknet_2_3_0_clock clknet_3_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_152_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _03882_ _05151_ _05164_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05603__A1 _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05603__B2 _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ _05113_ _05116_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09345__A2 _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08856__A1 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06331__A2 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05410_ _00847_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08608__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ _01648_ _01688_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08608__B2 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05341_ _00825_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05517__S1 _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08060_ _03261_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05272_ _00769_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_162_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07011_ mem.mem_dff.code_mem\[13\]\[0\] _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05842__A1 _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05842__B2 _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07993__I _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08387__A3 _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08962_ _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10843__CLK clknet_leaf_190_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07913_ _03132_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09336__A2 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08893_ _03973_ _03971_ _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_190_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07844_ _03090_ _03087_ _03082_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07942__B _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _02978_ _03032_ _03028_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10993__CLK clknet_leaf_13_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ _04281_ _04475_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06726_ _02201_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08329__I _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__B2 stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07233__I _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08311__A3 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09445_ net155 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06657_ mem.mem_dff.code_mem\[3\]\[6\] _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05889__S _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05608_ _01103_ _01154_ _01155_ _01134_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09376_ _01765_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06588_ _02102_ _02103_ _02092_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05530__B1 stack\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10406__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ mem.mem_dff.code_mem\[8\]\[6\] _03292_ _03293_ mem.mem_dff.code_mem\[22\]\[6\]
+ _03516_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_166_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05539_ _01087_ stack\[11\]\[6\] _01080_ stack\[10\]\[6\] _01040_ _01088_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10406__B2 stack\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08075__A2 _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09272__A1 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05688__I _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03450_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _02594_ _02590_ _02595_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05833__A1 _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05833__B2 _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08189_ mem.mem_dff.data_mem\[0\]\[1\] _03318_ _03319_ _03383_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _05059_ _05055_ _05060_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _04976_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05597__B1 stack\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05356__C _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06010__A1 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06010__B2 _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08239__I _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _00576_ clknet_4_3_0_clock net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10716__CLK clknet_leaf_36_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09263__A1 _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06077__A1 _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05824__A1 _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10009__I _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09015__A1 _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09015__B2 _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__CLK clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09566__A2 _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _00010_ clknet_leaf_39_clock mem.mem_dff.cycles\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _03858_ _04209_ _03189_ _03690_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_174_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07318__I mem.mem_dff.code_mem\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05978__I2 stack\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06222__I _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10333__B1 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05890_ _01280_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05282__B _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ mem.mem_dff.code_mem\[27\]\[7\] _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08149__I _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08829__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08829__B2 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _02040_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07491_ _02814_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _04177_ _04217_ _04226_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06442_ _01379_ _01397_ _01225_ _01975_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09161_ _03716_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09254__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06373_ _01905_ _01910_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08112_ mem.mem_dff.code_mem\[5\]\[0\] _02199_ _02649_ mem.mem_dff.code_mem\[20\]\[0\]
+ _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_175_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06068__A1 _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05324_ _00877_ net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09092_ _01824_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05301__I _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08043_ _02345_ net188 _01174_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__A1 _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05255_ _00809_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09006__B2 stack\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _04866_ _01878_ _04874_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07228__I mem.mem_dff.code_mem\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11021__CLK clknet_leaf_16_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ _04013_ _03995_ _04009_ stack\[13\]\[5\] _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _01892_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input22_I i_wb_addr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _03076_ _03072_ _03077_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _03023_ _03020_ _03024_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08059__I _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ _02169_ _02200_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10739__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _02968_ _02960_ _02969_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__A1 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07898__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04395_ _04365_ _04398_ _04400_ _04401_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _01723_ _01628_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_139_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10889__CLK clknet_leaf_181_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__B2 _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A3 _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05211__I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05806__A1 _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07847__B _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10203_ _04185_ _05045_ _05046_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_134_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11183_ net233 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06231__A1 _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _01216_ _04969_ _04973_ _04994_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _04922_ _04932_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05814__C _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08287__A2 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _00559_ clknet_leaf_129_clock net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06298__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10898_ _00490_ clknet_leaf_185_clock stack\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_173_clock_I clknet_4_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__A1 _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07798__A1 _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07757__B _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09528__I delay_cycles\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11044__CLK clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05992__S _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ mem.mem_dff.code_mem\[12\]\[3\] _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _03731_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05942_ _00900_ stack\[21\]\[4\] _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__B1 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09711__A2 _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _01892_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05873_ _00809_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _02824_ _02905_ _02898_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05959__S1 _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ stack\[31\]\[7\] _03727_ _03738_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07543_ mem.mem_dff.code_mem\[27\]\[3\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_207_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07474_ _02790_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07511__I _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ stack\[21\]\[0\] _04213_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06425_ _01649_ _01956_ _01961_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09227__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09144_ _03186_ _04025_ _04026_ _03691_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06356_ net13 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05307_ _00798_ _00858_ _00860_ _00816_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09242__A4 _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ _04040_ _04093_ _04096_ stack\[23\]\[6\] _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_175_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06287_ _01814_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08026_ _03230_ _03231_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05238_ _00784_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05895__S0 _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10411__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ _04857_ _04863_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07961__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06797__I _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08928_ _03898_ _04001_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09702__A2 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output226_I net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10561__CLK clknet_leaf_96_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08859_ _03781_ _03946_ _03948_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07713__A1 _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_6_0_clock clknet_3_3_0_clock clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _00413_ clknet_leaf_160_clock stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08269__A2 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10752_ _00344_ clknet_leaf_38_clock mem.io_data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _00275_ clknet_leaf_60_clock mem.mem_dff.data_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05342__I3 stack\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11067__CLK clknet_opt_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06452__A1 _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06204__B2 _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06755__A2 _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10904__CLK clknet_leaf_180_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05802__I1 stack\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _01215_ _04935_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ _00689_ clknet_leaf_6_clock net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09083__I _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06500__I _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10048_ net38 net39 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09457__A1 _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout257_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10178__B _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__I1 stack\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05333__I3 stack\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05987__S _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06210_ _01742_ _01743_ _01747_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05494__A2 stack\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07190_ mem.mem_dff.code_mem\[17\]\[6\] _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__CLK clknet_leaf_75_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05786__I _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06443__A1 _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06072_ _01607_ _01615_ _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06994__A2 _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09900_ _04598_ _04808_ _03183_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09831_ _04600_ _04762_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10584__CLK clknet_leaf_86_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__A1 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06974_ mem.mem_dff.code_mem\[12\]\[0\] _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09762_ exec.memory_input\[1\] _04286_ _04712_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07506__I _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ _03819_ _03826_ _03834_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05925_ stack\[14\]\[3\] stack\[15\]\[3\] _00770_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09693_ _01630_ _04258_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09696__A1 _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ _03781_ _03778_ _03773_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05856_ _01398_ _01399_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _03227_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09448__A1 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05787_ stack\[28\]\[0\] stack\[29\]\[0\] _01330_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07526_ _02755_ _02832_ _02842_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05309__I0 stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09999__A2 _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _02788_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08671__A2 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05897__S _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06408_ _01905_ _01941_ _01944_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_07388_ _02729_ _02733_ _02735_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09127_ _04122_ _04147_ _04149_ stack\[18\]\[1\] _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06339_ _01866_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09168__I _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06434__A1 _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08072__I _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ _03869_ _04095_ _04097_ _04098_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06434__B2 _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output176_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__CLK clknet_leaf_148_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ _03218_ _03209_ _03205_ stack\[28\]\[2\] _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10107__I _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11020_ _00612_ clknet_leaf_16_clock cycles_per_ms\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__A4 _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__B1 _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06320__I _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09687__A1 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05712__A3 _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05563__I3 stack\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10049__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10804_ _00396_ clknet_leaf_171_clock stack\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _00327_ clknet_leaf_64_clock mem.mem_dff.data_mem\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08662__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__CLK clknet_leaf_70_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10666_ _00258_ clknet_leaf_57_clock mem.mem_dff.code_mem\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _00189_ clknet_leaf_99_clock mem.mem_dff.code_mem\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06425__A1 _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05539__C _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11149_ _00741_ clknet_leaf_138_clock stack\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05787__I0 stack\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09127__B1 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__I _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09678__A1 _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05710_ _01232_ _01253_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06690_ _02174_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05641_ net131 _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08360_ mem.mem_dff.code_mem\[12\]\[7\] _02415_ _03432_ mem.mem_dff.code_mem\[14\]\[7\]
+ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08157__I _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05572_ _00979_ _01101_ _01111_ _01120_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ _02198_ _02586_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08291_ _03335_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07456__A3 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07242_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05467__A2 _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _02506_ _02565_ _02558_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09602__A1 _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01661_ _01666_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06416__A1 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06055_ _01144_ _01591_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09905__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09814_ _04413_ _04666_ _01125_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09745_ _04690_ _04702_ _04675_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ mem.mem_dff.code_mem\[11\]\[4\] _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05908_ stack\[22\]\[3\] stack\[23\]\[3\] _01403_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10279__A2 _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _04625_ _04626_ _04627_ _04635_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06888_ mem.mem_dff.code_mem\[9\]\[7\] _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__A1 _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05839_ _01010_ _01381_ _01382_ _01285_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08627_ _01932_ _03664_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05950__I0 stack\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08558_ _01763_ _03700_ _03705_ _03709_ _03710_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_208_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ mem.mem_dff.code_mem\[26\]\[4\] _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08489_ _01829_ _03632_ _03655_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09841__A1 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A2 _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06655__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10520_ _00112_ clknet_leaf_112_clock mem.mem_dff.code_mem\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05458__A2 _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10451_ _00043_ clknet_leaf_73_clock mem.mem_dff.code_mem\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06407__A1 _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__A2 _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10382_ _03215_ _05172_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11105__CLK clknet_leaf_35_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05630__A2 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11003_ _00595_ clknet_leaf_128_clock exec.memory_input\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08580__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05394__A1 _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08332__B2 mem.mem_dff.code_mem\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3_0_clock clknet_2_1_0_clock clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A2 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A1 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09832__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A2 _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06934__B _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _00310_ clknet_leaf_36_clock mem.mem_dff.data_mem\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__I _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _00241_ clknet_leaf_116_clock mem.mem_dff.code_mem\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08399__A1 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07071__A1 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09348__B1 _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10191__B _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _03102_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08166__A4 _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06811_ _02278_ _02273_ _02280_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07791_ _02963_ _03047_ _03039_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06742_ _02225_ _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09530_ delay_cycles\[6\] delay_cycles\[5\] delay_cycles\[4\] _04489_ _04490_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_114_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06895__I _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10622__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08323__B2 mem.mem_dff.code_mem\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ net157 _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06673_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05732__C _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10130__A1 _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08874__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10130__B2 _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ net125 _03588_ _03589_ _03090_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05624_ mem.select _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10210__I _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09392_ _04368_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08343_ mem.mem_dff.data_mem\[2\]\[6\] _03327_ _03375_ mem.mem_dff.data_mem\[6\]\[6\]
+ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10772__CLK clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05555_ _01077_ stack\[28\]\[6\] stack\[29\]\[6\] _01078_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09823__A1 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06844__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08274_ mem.mem_dff.code_mem\[19\]\[4\] _03366_ _03359_ mem.mem_dff.code_mem\[21\]\[4\]
+ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05486_ _00932_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08615__I _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06101__A3 _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07225_ _02370_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11128__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ mem.mem_dff.code_mem\[16\]\[6\] _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06107_ _01587_ _01650_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07087_ _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07601__A3 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05999__I0 stack\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input52_I i_wb_data[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09446__I _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06038_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A1 _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output139_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07989_ _03199_ _03200_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_216_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _04686_ _04676_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08314__B2 _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09659_ _04539_ _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10121__A1 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08865__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05679__A2 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05214__I _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__A3 _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09814__A1 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__A2 _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06754__B _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _00095_ clknet_leaf_107_clock mem.mem_dff.code_mem\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10434_ _00026_ clknet_leaf_75_clock mem.mem_dff.code_mem\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10188__A1 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09042__A2 _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__B1 _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _01923_ _05153_ _05161_ stack\[17\]\[5\] _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09356__I _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ _04191_ _05114_ _05115_ _04167_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10645__CLK clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06929__B _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07604__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10112__A1 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10795__CLK clknet_leaf_5_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08856__A2 _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10112__B2 _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05914__I0 stack\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09805__A1 _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08608__A2 _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05340_ _00892_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10186__B _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07292__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05271_ _00797_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07010_ _02435_ _02428_ _02438_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05995__S _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_170_clock clknet_4_3_0_clock clknet_leaf_170_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10179__A1 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09033__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__A1 _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09266__I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08170__I _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08961_ _03186_ _04025_ _04026_ _03234_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_185_clock clknet_4_4_0_clock clknet_leaf_185_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07912_ _03132_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08892_ _01715_ _03823_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_168_clock_I clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _02055_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10351__A1 _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ mem.mem_dff.data_mem\[1\]\[6\] _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _04474_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06725_ _02201_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08847__A2 _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06656_ _02157_ _02154_ _02158_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09444_ _04410_ _04416_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08311__A4 _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05905__I0 stack\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_123_clock clknet_4_12_0_clock clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ stack\[22\]\[7\] _01080_ _01076_ stack\[23\]\[7\] _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06587_ _02099_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09375_ _03242_ _04351_ _04352_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05530__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05530__B2 _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ _03513_ _03514_ _03515_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05538_ _00932_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10406__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10518__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08257_ mem.dff_data_out\[3\] _03449_ _03336_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05469_ _00937_ _01019_ _00879_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_clock clknet_4_7_0_clock clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07208_ _02506_ _02592_ _02583_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05833__A2 _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08188_ _03376_ _03380_ _03382_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07139_ _02506_ _02539_ _02528_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05918__B _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10668__CLK clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10150_ net163 _04999_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05597__A1 _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05597__B2 _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10081_ _04936_ _04948_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A1 _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _00575_ clknet_leaf_9_clock net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05521__A1 _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A2 _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08191__S _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09015__A2 _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10417_ _00009_ clknet_leaf_39_clock mem.mem_dff.cycles\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08774__A1 _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09971__B1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10348_ _05151_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05588__A1 _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _01888_ _05089_ _05101_ stack\[30\]\[4\] _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08526__A1 _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10333__A1 _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__B2 stack\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_clock clknet_4_8_0_clock clknet_leaf_40_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08829__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10097__B1 _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06510_ net244 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07490_ _02760_ _02813_ _02096_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_34_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0_0_clock clknet_0_clock clknet_2_0_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06441_ _01168_ _01968_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ _04173_ _04171_ _04174_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_55_clock clknet_4_12_0_clock clknet_leaf_55_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06372_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09254__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08111_ _03306_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06068__A2 _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05323_ _00876_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_94_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09091_ _04050_ _04115_ _04123_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05254_ _00785_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09006__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09993_ _02051_ _04867_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05457__C _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__CLK clknet_leaf_142_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07953__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08944_ _01922_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _03959_ _03942_ _03960_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09190__A1 _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _02963_ _03074_ _03066_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I i_la_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ _02963_ _03021_ _03011_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06708_ _02199_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _02952_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09493__A2 _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04374_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06639_ _02142_ _02139_ _02145_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _01214_ _04315_ _04335_ _04337_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ mem.mem_dff.code_mem\[19\]\[5\] _03366_ _03359_ mem.mem_dff.code_mem\[21\]\[5\]
+ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07256__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ _03241_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_2_0_clock clknet_3_1_0_clock clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07419__I _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _03202_ _03990_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11182_ net235 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06323__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10133_ _01169_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06231__A2 _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08508__A1 _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10064_ _04931_ _04920_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10315__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05990__A1 _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09181__A1 stack\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__B1 _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10966_ _00558_ clknet_leaf_129_clock net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09484__A2 _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10897_ _00489_ clknet_leaf_182_clock stack\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_116_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__I _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05353__S0 _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10983__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__A1 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06990_ _02422_ _02417_ _02423_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I i_la_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05941_ _01014_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09172__A1 _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09172__B2 stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05872_ _01302_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08660_ _03791_ _03774_ _03793_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09711__A3 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08514__A4 _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07611_ mem.mem_dff.code_mem\[29\]\[2\] _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05733__A1 _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _03737_ _03717_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07542_ _02854_ _02848_ _02855_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09475__A2 _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A1 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ mem.mem_dff.code_mem\[25\]\[4\] _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08683__B1 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09212_ _04212_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06424_ _01649_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A2 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ _03936_ _04157_ _04160_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06355_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07948__B _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08986__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05306_ _00783_ _00797_ _00859_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_09074_ _03663_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06286_ _01797_ _01642_ _01826_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05237_ _00791_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08025_ _01677_ _01925_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__S1 _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06213__A2 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09976_ delay_cycles\[22\] _04810_ _04859_ _04862_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08927_ _03995_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10706__CLK clknet_leaf_29_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09163__A1 _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _01639_ _03940_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__A2 _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08910__A1 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output121_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07809_ _02978_ _03058_ _03054_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05724__A1 _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output219_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _03893_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10820_ _00412_ clknet_leaf_170_clock stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10856__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _00343_ clknet_leaf_38_clock mem.io_data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10682_ _00274_ clknet_leaf_54_clock mem.mem_dff.data_mem\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07229__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08977__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10233__B1 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06452__A2 _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08729__A1 _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06053__I _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05412__B1 stack\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _04975_ _04141_ _04979_ _04980_ _04776_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_212_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_clock_I clknet_4_9_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11096_ _00688_ clknet_leaf_6_clock net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09154__A1 _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10047_ _00842_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08901__A1 _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08708__I _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__C _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10949_ _00541_ clknet_leaf_192_clock stack\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08968__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06140_ _01678_ _01680_ _01682_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09090__B1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10194__B _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07640__A1 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10729__CLK clknet_leaf_64_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09393__A1 exec.out_of_order_exec vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _04756_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07943__A2 _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09761_ _04713_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06973_ _02406_ _02398_ _02409_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09145__A1 _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08712_ _03776_ _03830_ _03833_ stack\[8\]\[0\] _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05924_ stack\[12\]\[3\] stack\[13\]\[3\] _01410_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09692_ _04650_ _04651_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10879__CLK clknet_leaf_143_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09696__A2 _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05855_ stack\[18\]\[6\] stack\[19\]\[6\] stack\[16\]\[6\] stack\[17\]\[6\] _00868_
+ _00890_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__05706__A1 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06847__B _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _03720_ _03706_ _03723_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_187_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05786_ _01329_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07525_ _02841_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05309__I1 stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07456_ _02787_ _02440_ _02069_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_211_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06407_ _01878_ _01871_ _01910_ _01943_ _01874_ _01873_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_202_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07387_ _02704_ _02734_ _02727_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input82_I rambus_wb_dat_i[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09126_ _04066_ _04144_ _04150_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01026_ _01811_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07631__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09057_ _03752_ _04092_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06269_ _00916_ _01809_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output169_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06198__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07934__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09959_ _04819_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05796__I1 stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09136__B2 stack\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10123__I _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09687__A2 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__B1 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06370__A1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11034__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10803_ _00395_ clknet_leaf_166_clock stack\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10049__A3 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _00326_ clknet_leaf_50_clock mem.mem_dff.data_mem\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08464__S _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ _00257_ clknet_leaf_77_clock mem.mem_dff.code_mem\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _00188_ clknet_leaf_99_clock mem.mem_dff.code_mem\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06425__A2 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05633__B1 intr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08178__A2 _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07925__A2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06511__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _00740_ clknet_leaf_138_clock stack\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09127__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__B2 stack\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11079_ _00671_ clknet_leaf_125_clock delay_counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07689__A1 _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__B1 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05640_ net132 _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05571_ _00950_ _01119_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07310_ mem.mem_dff.code_mem\[21\]\[0\] _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ _03474_ _03481_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06113__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07241_ _02532_ _02620_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07861__A1 _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ mem.mem_dff.code_mem\[17\]\[1\] _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08173__I _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10551__CLK clknet_leaf_79_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _01662_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_145_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__A1 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ net189 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05778__I1 _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09744_ _04678_ _04701_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06956_ _02393_ _02385_ _02396_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05907_ stack\[20\]\[3\] stack\[21\]\[3\] _00791_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09675_ _04571_ _04634_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08877__B1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06887_ _02339_ _02334_ _02340_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08626_ _03765_ _03766_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05838_ stack\[8\]\[7\] stack\[9\]\[7\] _00800_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10099__B _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08557_ _03215_ _03707_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05769_ _01258_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05950__I1 stack\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07508_ _02826_ _02817_ _02828_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ _03654_ _03642_ _03648_ stack\[19\]\[3\] _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09841__A2 _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A3 _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ _02763_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _00042_ clknet_leaf_69_clock mem.mem_dff.code_mem\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08083__I _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _04133_ _04134_ _04136_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10381_ stack\[15\]\[1\] _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09907__I _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11002_ _00594_ clknet_leaf_127_clock exec.memory_input\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_2_0_clock_I clknet_3_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05918__A1 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09109__A1 _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06591__A1 _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05394__A2 _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08868__B1 _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08332__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10424__CLK clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__A1 _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06343__B2 _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10574__CLK clknet_leaf_89_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10717_ _00309_ clknet_leaf_36_clock mem.mem_dff.data_mem\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09089__I _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06506__I _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10648_ _00240_ clknet_leaf_116_clock mem.mem_dff.code_mem\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05410__I _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08399__A2 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10579_ _00171_ clknet_leaf_84_clock mem.mem_dff.code_mem\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06950__B _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09817__I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05606__B1 stack\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__A1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__B2 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05909__A1 _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05909__B2 _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06810_ _02279_ _02274_ _02270_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07790_ mem.mem_dff.data_mem\[2\]\[1\] _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06741_ _02095_ _02224_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09460_ _04428_ _04430_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06672_ _02095_ _02171_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06334__A1 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10130__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08411_ _03568_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05623_ _01170_ net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09391_ _04367_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10917__CLK clknet_leaf_147_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ mem.mem_dff.code_mem\[0\]\[6\] _03451_ _03523_ _03531_ _03473_ _03532_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05554_ _01041_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08273_ mem.mem_dff.code_mem\[2\]\[4\] _03349_ _03350_ mem.mem_dff.code_mem\[18\]\[4\]
+ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07834__A1 _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05485_ _01033_ _01034_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ mem.mem_dff.code_mem\[18\]\[5\] _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06101__A4 _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__B1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _02552_ _02549_ _02553_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06106_ _01596_ _01603_ _01614_ _01620_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_07086_ _02287_ _02412_ _02255_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05999__I1 stack\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06037_ _01231_ _01253_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07247__I _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input45_I i_wb_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A2 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10447__CLK clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _01633_ _01635_ _01604_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_210_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_89_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _04685_ _04257_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06939_ _02382_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09658_ _04550_ _04548_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10121__A2 _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10597__CLK clknet_leaf_99_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output201_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ _03751_ _03753_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05679__A3 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09589_ _04540_ _04541_ _04548_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08078__A1 _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__I _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09814__A2 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06628__A2 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10502_ _00094_ clknet_leaf_108_clock mem.mem_dff.code_mem\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09027__B1 _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05230__I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10433_ _00025_ clknet_leaf_76_clock mem.mem_dff.code_mem\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__I _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _03879_ _05151_ _05163_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08250__B2 _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10295_ _05110_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08305__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08856__A3 _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05914__I1 stack\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07620__I _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05270_ _00783_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__B _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10179__A2 _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08241__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06252__B1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08960_ _01691_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07911_ mem.mem_dff.data_mem\[5\]\[4\] _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _03780_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ mem.mem_dff.data_mem\[3\]\[5\] _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_90_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10351__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07773_ _03034_ _03031_ _03035_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09512_ _04323_ _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06724_ mem.mem_dff.code_mem\[5\]\[4\] _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10221__I _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06307__A1 exec.memory_input\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04406_ _04415_ _02000_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06655_ _02122_ _02155_ _02151_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__B _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05905__I1 stack\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05606_ _01077_ stack\[20\]\[7\] stack\[21\]\[7\] _01078_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ mem.io_data_out\[7\] _04320_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09257__B1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06586_ _02101_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07530__I _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05530__A2 stack\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ mem.mem_dff.code_mem\[23\]\[6\] _03391_ _03392_ mem.mem_dff.code_mem\[31\]\[6\]
+ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05537_ _01062_ _01085_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08256_ _03443_ _03448_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09009__B1 _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06146__I _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05468_ stack\[27\]\[4\] stack\[24\]\[4\] stack\[25\]\[4\] stack\[26\]\[4\] _00953_
+ _00954_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08480__A1 _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ mem.mem_dff.code_mem\[18\]\[1\] _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08187_ mem.mem_dff.data_mem\[4\]\[1\] _03101_ _03131_ mem.mem_dff.data_mem\[5\]\[1\]
+ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05399_ stack\[11\]\[3\] stack\[8\]\[3\] stack\[9\]\[3\] stack\[10\]\[3\] _00942_
+ _00928_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07138_ mem.mem_dff.code_mem\[16\]\[1\] _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08232__A1 mem.mem_dff.code_mem\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07035__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07069_ _02365_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05841__I0 stack\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10080_ _04921_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09732__A1 _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06546__A1 _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__A2 _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10982_ _00574_ clknet_leaf_9_clock net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__I _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09248__B1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08536__I _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10612__CLK clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _00008_ clknet_leaf_40_clock mem.dff_data_ready vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07026__A2 _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08774__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _03668_ _01637_ _03630_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_112_clock_I clknet_4_12_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10278_ _05059_ _05098_ _05102_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10762__CLK clknet_leaf_49_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08526__A2 _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10333__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07615__I _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11118__CLK clknet_leaf_141_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10097__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10097__B2 intr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05899__I0 stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06440_ _01937_ _01974_ _01749_ _01975_ _01816_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10197__B _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06371_ _01842_ _01906_ _01908_ _01902_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08110_ mem.mem_dff.code_mem\[1\]\[0\] _02070_ _02561_ mem.mem_dff.code_mem\[17\]\[0\]
+ _02026_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_37_clock_I clknet_4_11_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05322_ _00875_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09090_ _04122_ _04117_ _04120_ stack\[24\]\[1\] _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ net253 _03243_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05253_ _00799_ _00804_ _00807_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08214__A1 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05418__I3 stack\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09992_ _02998_ _04869_ _04873_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06776__A1 _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _03959_ _04003_ _04012_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08874_ _03842_ _03946_ _03955_ stack\[26\]\[4\] _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07525__I _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10324__A2 _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07825_ mem.mem_dff.data_mem\[3\]\[1\] _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09190__A2 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ mem.mem_dff.data_mem\[1\]\[1\] _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06707_ _02025_ _02198_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07687_ _02044_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ _04313_ _04399_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06638_ _02144_ _02140_ _02130_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ _04336_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06569_ _02056_ _02085_ _02081_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08308_ mem.mem_dff.code_mem\[2\]\[5\] _03349_ _03350_ mem.mem_dff.code_mem\[18\]\[5\]
+ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10635__CLK clknet_leaf_100_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__S _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08453__A1 _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _04268_ mem.dff_data_out\[0\] _04272_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output199_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10260__A1 _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ _02468_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09187__I _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10785__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _03635_ _03701_ _03994_ _03192_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11181_ net237 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09915__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ net157 _04961_ _04986_ _04572_ _04140_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08508__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ net36 net38 net39 _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07435__I _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10315__A2 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09181__A2 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09650__I cycles_per_ms\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10079__A1 _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10079__B2 intr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10965_ _00557_ clknet_leaf_192_clock stack\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08692__A1 _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10896_ _00488_ clknet_leaf_180_clock stack\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_184_clock clknet_4_4_0_clock clknet_leaf_184_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_197_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08444__A1 _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10251__A1 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05353__S1 _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10003__A1 _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06758__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_122_clock clknet_4_9_0_clock clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _01259_ _01483_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10306__A2 _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09172__A2 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10508__CLK clknet_leaf_108_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05871_ _01409_ _01411_ _01413_ _01414_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09711__A4 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07610_ _02907_ _02904_ _02908_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_208_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08590_ _01975_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05733__A2 _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07541_ _02824_ _02849_ _02842_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07472_ _02798_ _02791_ _02800_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08683__A1 _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08683__B2 stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09211_ _04185_ _04210_ _04211_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05497__A1 _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06423_ _01959_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ _03937_ _04142_ _04153_ stack\[18\]\[7\] _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08435__A1 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06354_ _01891_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05305_ stack\[27\]\[1\] stack\[24\]\[1\] stack\[25\]\[1\] stack\[26\]\[1\] _00856_
+ _00793_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08986__A2 _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09073_ _03230_ _03661_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06285_ stack\[2\]\[2\] _01718_ _01825_ _01759_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_200_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08024_ _01692_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05236_ _00790_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07964__B _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09975_ _04501_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08926_ stack\[13\]\[0\] _03999_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07255__I _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09163__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08857_ _03946_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__B1 _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07808_ mem.mem_dff.data_mem\[2\]\[6\] _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08910__A2 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ _01639_ _03807_ _02008_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_166_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05724__A2 stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ _03007_ _03002_ _03008_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output114_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10750_ _00342_ clknet_leaf_38_clock mem.io_data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08674__A1 stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05503__I _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _03624_ _04384_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ _00273_ clknet_leaf_51_clock mem.mem_dff.data_mem\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08426__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10233__A1 _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08977__A2 _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10233__B2 stack\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__A2 _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05412__A1 _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05412__B2 _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10115_ _04103_ _04973_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11095_ _00687_ clknet_leaf_6_clock net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_clock clknet_4_12_0_clock clknet_leaf_54_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10046_ _04888_ _04913_ _04914_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07165__A1 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__A2 _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10800__CLK clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_clock clknet_4_14_0_clock clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08114__B1 _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10948_ _00540_ clknet_leaf_192_clock stack\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__A1 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10879_ _00471_ clknet_leaf_143_clock stack\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08417__A1 _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10224__A1 _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08968__A2 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09090__A1 _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09090__B2 stack\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _01608_ _01609_ _01611_ _01613_ _01582_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA_clkbuf_0_clock_I clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ exec.memory_input\[0\] _04276_ _04712_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06972_ _02407_ _02399_ _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08711_ _03832_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09145__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05923_ _01302_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09691_ delay_counter\[0\] delay_counter\[1\] delay_counter\[3\] delay_counter\[2\]
+ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_187_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08642_ _01643_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10480__CLK clknet_leaf_123_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05854_ _01258_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ _03224_ _03711_ _03722_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05785_ _00899_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08105__B1 _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07524_ _02840_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08656__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05309__I2 stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05323__I _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ _02022_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06406_ _01872_ _01942_ _01909_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_210_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07386_ _02732_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ _04024_ _04147_ _04149_ stack\[18\]\[0\] _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06337_ _01872_ _01875_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_176_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input75_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ stack\[23\]\[1\] _04096_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06268_ _01732_ _01634_ _01734_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08007_ _01823_ _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05219_ net137 _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06199_ _01740_ _01741_ _01730_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_clock_I clknet_2_1_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_6_clock_I clknet_4_2_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09958_ _04850_ _04851_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05945__A2 stack\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_159_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10823__CLK clknet_leaf_160_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09136__A2 _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ stack\[10\]\[6\] _03976_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09889_ _04500_ _04768_ _04795_ net57 _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08344__B1 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__A1 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08895__B2 stack\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10973__CLK clknet_leaf_43_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10802_ _00394_ clknet_leaf_167_clock stack\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08647__A1 _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10049__A4 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10733_ _00325_ clknet_leaf_49_clock mem.mem_dff.data_mem\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10664_ _00256_ clknet_leaf_77_clock mem.mem_dff.code_mem\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08544__I _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05881__A1 _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09072__A1 _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10595_ _00187_ clknet_leaf_99_clock mem.mem_dff.code_mem\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08178__A3 _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11147_ _00739_ clknet_leaf_191_clock stack\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05408__I _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__A2 _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11078_ _00670_ clknet_leaf_132_clock delay_counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10029_ _04898_ _04900_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__A1 _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07623__I mem.mem_dff.code_mem\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__B2 _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05570_ _01102_ _01112_ _01116_ _01118_ _01089_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07779__B _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06683__B _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06113__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ _02619_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07171_ _02560_ _02564_ _02566_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__A1 stack\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06122_ _01663_ _01664_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_199_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__A1 _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ _01596_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__I mem.sram_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10846__CLK clknet_leaf_161_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09366__A2 _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09812_ _01173_ _04744_ _04748_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07019__B _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_160_clock_I clknet_4_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05927__A2 _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06955_ _02394_ _02386_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09743_ _04691_ _04700_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07129__A1 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10996__CLK clknet_leaf_8_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05906_ _01398_ _01449_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09674_ _04578_ _04633_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06886_ _02279_ _02335_ _02331_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08877__A1 _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__B2 stack\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ net149 _03763_ _03760_ stack\[3\]\[5\] _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08341__A3 _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05837_ stack\[10\]\[7\] stack\[11\]\[7\] _00868_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06149__I _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__A1 _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08556_ stack\[31\]\[1\] _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05768_ _01310_ _01311_ _00944_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05560__B1 _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07507_ _02742_ _02819_ _02827_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _03220_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05699_ _01206_ _01199_ _01242_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07438_ mem.mem_dff.code_mem\[24\]\[4\] _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05863__A1 _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_85_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07369_ mem.mem_dff.code_mem\[22\]\[5\] _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09054__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _04135_ _04118_ _04127_ stack\[24\]\[6\] _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_202_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output181_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08801__A1 _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _01352_ _05171_ _05173_ _05175_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05615__A1 _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09039_ _04040_ _04072_ _04078_ stack\[9\]\[6\] _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05615__B2 stack\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07708__I _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11001_ _00593_ clknet_leaf_128_clock exec.memory_input\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05228__I _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__A1 _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__B2 _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11001__CLK clknet_leaf_128_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_6_0_clock_I clknet_3_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08868__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__B2 stack\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11151__CLK clknet_4_7_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__A3 _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10719__CLK clknet_leaf_30_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09293__A1 _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05898__I _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10716_ _00308_ clknet_leaf_36_clock mem.mem_dff.data_mem\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10647_ _00239_ clknet_leaf_116_clock mem.mem_dff.code_mem\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10578_ _00170_ clknet_leaf_89_clock mem.mem_dff.code_mem\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05606__A1 _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05606__B2 _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07618__I mem.mem_dff.code_mem\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A2 _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06522__I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10363__B1 _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06740_ _02170_ net229 _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08449__I _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_4_1_clock clknet_opt_4_0_clock clknet_opt_4_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09520__A2 _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06671_ _02170_ net227 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08410_ _03581_ _03590_ _03593_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05622_ _01169_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _01198_ _01200_ _01202_ _01575_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05542__B1 stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05802__S _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _03524_ _03529_ _03530_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05553_ _01028_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09284__A1 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__B2 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ mem.mem_dff.code_mem\[5\]\[4\] _03352_ _03353_ mem.mem_dff.code_mem\[20\]\[4\]
+ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08184__I _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05484_ _01030_ stack\[16\]\[5\] stack\[17\]\[5\] _01031_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ _02602_ _02603_ _02606_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08117__C _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05845__A1 _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09036__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09036__B2 stack\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _02489_ _02550_ _02546_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08912__I _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07598__A1 _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06105_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07085_ mem.mem_dff.code_mem\[15\]\[0\] _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06036_ _01578_ _01579_ _01573_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11024__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10354__B1 _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06022__A1 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input38_I i_wb_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06022__B2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _01701_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06938_ _02288_ _02319_ _02381_ _02135_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09726_ _04250_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10106__B1 _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06869_ _02326_ _02323_ _02327_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09657_ _04529_ _04531_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06325__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08608_ _03752_ _03748_ _03749_ net145 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09588_ _04542_ _04543_ _04547_ cycles_per_ms\[12\] _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05679__A4 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _03694_ _03680_ _03687_ stack\[29\]\[6\] _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09275__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__I _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06628__A3 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10501_ _00093_ clknet_leaf_108_clock mem.mem_dff.code_mem\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09027__A1 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09027__B2 stack\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10432_ _00024_ clknet_leaf_76_clock mem.mem_dff.code_mem\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10363_ _01888_ _05153_ _05161_ stack\[17\]\[4\] _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10294_ _05109_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10345__B1 _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09750__A2 _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10541__CLK clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07513__A1 _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__A4 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10691__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06517__I _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09828__I _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11047__CLK clknet_leaf_26_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A2 _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07348__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__A1 stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06252__B2 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _03140_ _03133_ _03142_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08890_ _03971_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06004__A1 _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _03084_ _03085_ _03088_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_33_clock_I clknet_4_10_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09741__A2 _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ _02947_ _03032_ _03028_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06723_ _02209_ _02202_ _02211_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09511_ _03616_ _04437_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06307__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04411_ _04361_ _04414_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06654_ mem.mem_dff.code_mem\[3\]\[5\] _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05605_ _01129_ _01151_ _01152_ _01127_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09373_ _04283_ mem.dff_data_out\[7\] _04350_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06585_ net249 _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ mem.mem_dff.code_mem\[6\]\[6\] _03388_ _03389_ mem.mem_dff.code_mem\[30\]\[6\]
+ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05536_ _01083_ stack\[8\]\[6\] stack\[9\]\[6\] _01084_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06427__I _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08255_ mem.mem_dff.data_mem\[0\]\[3\] _03318_ _03319_ _03447_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09009__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05467_ stack\[30\]\[4\] _00925_ _00993_ stack\[31\]\[4\] _00961_ _01018_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__09009__B2 stack\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08480__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06871__B _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ _02585_ _02590_ _02593_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _02290_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08642__I _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05398_ _00781_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07137_ _02530_ _02538_ _02540_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10414__CLK clknet_4_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ _02470_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07991__A1 _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06019_ _01342_ _01559_ _01562_ _01480_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05841__I1 stack\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__B1 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09193__B1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09732__A2 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output144_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10564__CLK clknet_leaf_82_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06546__A2 _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _04353_ _04668_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_210_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10981_ _00573_ clknet_leaf_44_clock net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09496__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05506__B1 stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09248__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09248__B2 stack\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__A1 _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__C1 mem.mem_dff.code_mem\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08552__I _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10415_ _00007_ clknet_leaf_3_clock stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06234__A1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10346_ _03854_ _05148_ _05150_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10907__CLK clknet_leaf_186_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05832__I1 stack\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _01857_ _05090_ _05101_ stack\[30\]\[3\] _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_215_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05416__I _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__A1 _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09239__A1 _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05899__I1 stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06370_ _01840_ _01907_ _01073_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05321_ _00874_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__CLK clknet_leaf_73_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ _03243_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05276__A2 _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05252_ _00806_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08462__I _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10587__CLK clknet_leaf_81_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _04870_ _01835_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ _04011_ _03995_ _04009_ stack\[13\]\[4\] _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_174_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06710__I _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08873_ _01860_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07824_ _03068_ _03072_ _03075_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07755_ _03013_ _03020_ _03022_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__A1 _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06706_ _02170_ net228 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05339__I0 stack\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07686_ mem.mem_dff.code_mem\[31\]\[3\] _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06637_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09425_ _04363_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06157__I _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06568_ mem.mem_dff.code_mem\[1\]\[5\] _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09356_ _02003_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08307_ mem.mem_dff.code_mem\[5\]\[5\] _03352_ _03353_ mem.mem_dff.code_mem\[20\]\[5\]
+ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05519_ _01063_ _01066_ _01068_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09287_ _04269_ _04271_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06499_ _02030_ _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08453__A2 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ mem.mem_dff.code_mem\[7\]\[3\] _03428_ _03429_ mem.mem_dff.code_mem\[9\]\[3\]
+ mem.mem_dff.code_mem\[28\]\[3\] _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10260__A2 _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08169_ _02136_ _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09402__A1 exec.out_of_order_exec vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10200_ _05043_ _05044_ _02005_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11180_ net240 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _04990_ _04141_ _04991_ _04992_ _04776_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_171_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05945__B _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09166__B1 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06620__I _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _04923_ _04924_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09931__I _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05236__I _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__A1 _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06776__B _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__I _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _00556_ clknet_leaf_188_clock stack\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07451__I _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10895_ _00487_ clknet_leaf_148_clock stack\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08692__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__A1 _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10251__A2 _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10003__A2 _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07955__A1 mem.mem_dff.data_mem\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10329_ _05138_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07626__I mem.mem_dff.code_mem\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08904__B1 _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ _01285_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07540_ mem.mem_dff.code_mem\[27\]\[2\] _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08132__A1 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07471_ _02742_ _02792_ _02799_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09880__A1 _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10001__B _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__B2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09210_ _03996_ _04087_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06422_ _01721_ net63 _01958_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09141_ _03963_ _04157_ _04158_ _04159_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06353_ _01890_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05304_ stack\[31\]\[1\] stack\[28\]\[1\] stack\[29\]\[1\] stack\[30\]\[1\] _00857_
+ _00847_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__06446__A1 exec.memory_input\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _03882_ _04095_ _04107_ _04108_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06284_ _01824_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08023_ _01893_ _03212_ _03229_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05235_ net135 _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_200_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08199__A1 mem.mem_dff.code_mem\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08199__B2 mem.mem_dff.code_mem\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08920__I _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_2_0_clock_I clknet_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09974_ _04857_ _04861_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ _03998_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03672_ _03673_ _03944_ _03945_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_input20_I i_wb_addr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__B2 _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07807_ _03060_ _03057_ _03061_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05999_ stack\[18\]\[1\] stack\[19\]\[1\] stack\[16\]\[1\] stack\[17\]\[1\] _00827_
+ _00828_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08787_ _01677_ _01685_ _01930_ _01713_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06921__A2 _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10602__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07738_ mem.mem_dff.data_mem\[0\]\[6\] _03003_ _02999_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07271__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05980__I0 stack\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07669_ _02870_ _02944_ _02953_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08674__A2 _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09408_ _04364_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10680_ _00272_ clknet_leaf_51_clock mem.mem_dff.data_mem\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10752__CLK clknet_leaf_38_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ _03241_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10233__A2 _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07937__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11163_ _00755_ clknet_leaf_5_clock stack\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05412__A2 stack\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10114_ _01191_ _04935_ _04941_ edge_interrupts _04978_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11094_ _00686_ clknet_leaf_14_clock net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10045_ delay_counter\[7\] _04882_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08362__A1 mem.mem_dff.code_mem\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05971__I0 stack\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10947_ _00539_ clknet_leaf_182_clock stack\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09862__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08665__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _00470_ clknet_leaf_143_clock stack\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06428__A1 stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10224__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09090__A2 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10047__I _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05651__A2 _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09917__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07356__I _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06600__A1 _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06971_ _02377_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ _03781_ _03829_ _03831_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05922_ _01426_ _01464_ _01465_ _01430_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10625__CLK clknet_leaf_104_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09690_ delay_counter\[5\] delay_counter\[4\] delay_counter\[7\] delay_counter\[6\]
+ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__A1 mem.mem_dff.code_mem\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08353__B2 mem.mem_dff.code_mem\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05853_ _01387_ _01396_ _00777_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08641_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10160__A1 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05784_ _00941_ _01326_ _01327_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08572_ _03721_ _03717_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05962__I0 stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ _01997_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10775__CLK clknet_leaf_122_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08656__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05309__I3 stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07454_ mem.mem_dff.code_mem\[25\]\[0\] _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09520__B _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__I _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06405_ _01901_ _01908_ _01902_ _01906_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07385_ _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09124_ _04148_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06336_ _01873_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09055_ _04089_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06267_ _01784_ _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08006_ _01764_ _03213_ _03216_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05218_ net138 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input68_I i_wb_we vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__A2 _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06198_ _01738_ _01739_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__A1 stack\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06170__I _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09957_ delay_cycles\[15\] _04846_ _04843_ _04531_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_183_clock clknet_4_4_0_clock clknet_leaf_183_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ _01933_ _03849_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_6_0_clock_I clknet_2_3_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_81_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output224_I net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08839_ _03724_ _03919_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08895__A2 _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05514__I _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10801_ _00393_ clknet_leaf_163_clock stack\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09844__A1 _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08647__A2 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10732_ _00324_ clknet_leaf_49_clock mem.mem_dff.data_mem\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _00255_ clknet_leaf_77_clock mem.mem_dff.code_mem\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10594_ _00186_ clknet_leaf_90_clock mem.mem_dff.code_mem\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09072__A2 _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07083__A1 _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07885__B _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__I _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05633__A2 intr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11080__CLK clknet_leaf_125_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08178__A4 _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10648__CLK clknet_leaf_116_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11146_ _00738_ clknet_leaf_191_clock stack\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05397__A1 _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11077_ _00669_ clknet_leaf_132_clock delay_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09391__I _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08335__B2 mem.mem_dff.code_mem\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ delay_counter\[4\] _04649_ _04899_ _01027_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10142__A1 _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10798__CLK clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout255_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__A1 _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08735__I _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02472_ _02565_ _02558_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06255__I _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09063__A2 _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06121_ net37 net6 _01654_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06121__I0 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__A2 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06052_ _01589_ _01592_ _01594_ _01595_ _01581_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_173_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09811_ _04417_ _04740_ _04741_ _04747_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_154_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_103_clock_I clknet_4_13_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _01168_ _01969_ _04694_ _04699_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06954_ _02377_ _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07129__A2 _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05905_ stack\[18\]\[3\] stack\[19\]\[3\] stack\[16\]\[3\] stack\[17\]\[3\] _00800_
+ _00890_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09673_ _04608_ _04594_ _04605_ _04632_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06885_ mem.mem_dff.code_mem\[9\]\[6\] _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08877__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _03724_ _03748_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05836_ _01281_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05767_ _00926_ stack\[27\]\[2\] _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08555_ _01182_ _03700_ _03706_ _01326_ _03708_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__A1 _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__A2 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__B2 stack\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07506_ _02783_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _01797_ _03632_ _03653_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05698_ _01216_ _01217_ _01233_ _01185_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07437_ _02771_ _02764_ _02773_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_13_0_clock_I clknet_3_6_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_clock clknet_4_9_0_clock clknet_leaf_53_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07368_ _02715_ _02716_ _02719_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07065__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ _01124_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06319_ _01829_ _01642_ _01858_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ mem.mem_dff.code_mem\[20\]\[5\] _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08801__A2 _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05615__A2 stack\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08380__I _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _04015_ _03849_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output174_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05937__C _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68_clock clknet_4_14_0_clock clknet_leaf_68_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_219_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11000_ _00592_ clknet_leaf_128_clock exec.memory_input\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10372__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10940__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06040__A2 _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08317__A1 mem.mem_dff.data_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A1 _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__B2 _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__A2 _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09293__A2 _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10715_ _00307_ clknet_leaf_31_clock mem.mem_dff.data_mem\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10646_ _00238_ clknet_leaf_117_clock mem.mem_dff.code_mem\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10577_ _00169_ clknet_leaf_91_clock mem.mem_dff.code_mem\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10470__CLK clknet_leaf_57_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06803__A1 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05606__A2 stack\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__C _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__B1 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10325__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10363__A1 _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11129_ _00721_ clknet_leaf_173_clock stack\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08308__A1 mem.mem_dff.code_mem\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10115__A1 _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__A2 _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__I _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06670_ net255 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_149_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05621_ _01168_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A1 _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09808__A1 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05542__B2 _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08340_ mem.mem_dff.code_mem\[11\]\[6\] _03299_ _02415_ mem.mem_dff.code_mem\[12\]\[6\]
+ mem.mem_dff.code_mem\[26\]\[6\] _03300_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05552_ _01082_ _01090_ _01100_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08465__I _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _03462_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05483_ _00925_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08492__B1 _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07222_ _02604_ _02605_ _02600_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10813__CLK clknet_leaf_159_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ mem.mem_dff.code_mem\[16\]\[5\] _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08244__B1 _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08795__A1 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _01647_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ _02493_ _02484_ _02496_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06035_ _01322_ _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05329__I _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10354__A1 _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10354__B2 stack\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _03194_ _03195_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07544__I _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09725_ _04388_ _04473_ _04665_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06937_ _02133_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10106__A1 _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05781__A1 _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10106__B2 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05781__B2 _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _04539_ _04549_ _04553_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05908__I0 stack\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06868_ _02264_ _02324_ _02315_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08607_ _03214_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05819_ _00786_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09587_ _04532_ _04546_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05533__A1 _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06799_ _02268_ _02260_ _02271_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _03237_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _03638_ _01703_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10493__CLK clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _00092_ clknet_leaf_108_clock mem.mem_dff.code_mem\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09027__A2 _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _00023_ clknet_leaf_76_clock mem.mem_dff.code_mem\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _01828_ _05152_ _05162_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10293_ stack\[27\]\[0\] _05112_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05239__I _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10345__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07454__I mem.mem_dff.code_mem\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05772__A1 _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08710__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10836__CLK clknet_leaf_189_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__A1 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10281__B1 _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__A1 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10986__CLK clknet_leaf_9_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _00221_ clknet_leaf_102_clock mem.mem_dff.code_mem\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07629__I mem.mem_dff.code_mem\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06252__A2 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10336__A1 _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07201__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07840_ _03086_ _03087_ _03082_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07364__I _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ mem.mem_dff.data_mem\[1\]\[5\] _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09510_ _04469_ _04471_ _04472_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06722_ _02150_ _02203_ _02210_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09441_ _04413_ _04323_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06653_ _02153_ _02154_ _02156_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05604_ stack\[18\]\[7\] _01140_ _01141_ stack\[19\]\[7\] _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06708__I _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09372_ _04348_ _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06584_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09257__A2 _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07268__A1 _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ mem.mem_dff.code_mem\[15\]\[6\] _03368_ _03369_ mem.mem_dff.code_mem\[29\]\[6\]
+ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05535_ _01015_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10272__B1 _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08254_ _03444_ _03445_ _03446_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05466_ _01009_ _01016_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09009__A2 _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07205_ _02591_ _02592_ _02583_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05768__B _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08185_ mem.mem_dff.data_mem\[1\]\[1\] _03377_ _03378_ mem.mem_dff.data_mem\[3\]\[1\]
+ mem.mem_dff.data_mem\[7\]\[1\] _03379_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05397_ _00920_ _00936_ _00948_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07136_ _02472_ _02539_ _02528_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07067_ mem.mem_dff.code_mem\[14\]\[4\] _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input50_I i_wb_data[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11141__CLK clknet_leaf_138_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06018_ _01476_ _01560_ _01561_ _01394_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__07991__A2 _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A1 _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10327__B2 _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09193__B2 stack\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08940__A1 _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output137_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ _03007_ _03178_ _03182_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09708_ _04322_ _04333_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10980_ _00572_ clknet_leaf_44_clock net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10859__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09496__A2 _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _04598_ cycles_per_ms\[0\] _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05506__A1 _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05357__I1 stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05506__B2 _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06618__I _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09248__A2 _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05809__A2 stack\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__C2 _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_opt_4_0_clock clknet_4_10_0_clock clknet_opt_4_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10414_ _00006_ clknet_4_3_0_clock stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10345_ _04994_ _05138_ _05145_ stack\[16\]\[7\] _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__A1 stack\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10276_ _05094_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05993__A1 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05993__B2 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07912__I _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08695__B1 _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09239__A2 _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05432__I _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__CLK clknet_leaf_127_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06972__B _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09839__I _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05320_ _00862_ _00873_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10254__B1 _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05251_ _00805_ _00782_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_175_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__S _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09990_ _04866_ _01837_ _04872_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ _01887_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08872_ _03957_ _03943_ _03958_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07094__I _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__B _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07823_ _03073_ _03074_ _03066_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07754_ _02930_ _03021_ _03011_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06705_ mem.mem_dff.code_mem\[5\]\[0\] _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05770__C _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ _02965_ _02959_ _02966_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05339__I1 stack\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ _04369_ _04396_ _04397_ _04382_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06636_ net247 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06161__A1 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09355_ _04303_ _04333_ _04334_ _04301_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06567_ _02083_ _02084_ _02086_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08306_ mem.mem_dff.code_mem\[1\]\[5\] _02071_ _03405_ mem.mem_dff.code_mem\[16\]\[5\]
+ _02027_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10245__B1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08989__A1 stack\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I rambus_wb_dat_i[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05518_ _00938_ _01067_ _00974_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09286_ net85 _00761_ _00762_ net108 _04270_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_21_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ net249 _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07661__A1 _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08237_ _02875_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05449_ _00950_ _00992_ _00999_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_166_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ mem.mem_dff.code_mem\[6\]\[1\] _02226_ _02731_ mem.mem_dff.code_mem\[23\]\[1\]
+ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08205__A3 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07119_ _02521_ _02516_ _02524_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08099_ mem.mem_dff.code_mem\[15\]\[0\] _02499_ _02902_ mem.mem_dff.code_mem\[29\]\[0\]
+ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _01217_ _04969_ _04973_ _01125_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05945__C _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ net18 net29 _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09166__B2 stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10681__CLK clknet_leaf_51_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_151_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08913__A1 stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__C1 mem.mem_dff.data_mem\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09469__A2 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11037__CLK clknet_leaf_33_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10963_ _00555_ clknet_leaf_184_clock stack\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06348__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10894_ _00486_ clknet_leaf_148_clock stack\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_76_clock_I clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07179__I _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07404__A1 _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07907__I mem.mem_dff.data_mem\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09394__I _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10328_ _05136_ _05139_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08231__C _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A1 _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10259_ _04206_ _05076_ _05082_ stack\[14\]\[7\] _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__05427__I _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08904__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__B2 stack\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__I _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06391__A1 _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05590__C _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__B1 _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08132__A2 _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ _02783_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09880__A2 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06421_ _01723_ _01957_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07891__A1 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09140_ _03238_ _04142_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06352_ _01072_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09093__B1 _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05303_ _00856_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07643__A1 _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ stack\[23\]\[5\] _04090_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06283_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06446__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08840__B1 _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07089__I _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06207__B _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08022_ _03228_ _03193_ _03225_ stack\[28\]\[5\] _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05234_ _00788_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06721__I _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ delay_cycles\[21\] _04810_ _04859_ _04503_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05957__A1 _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09148__A1 stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08924_ _03973_ _03995_ _03997_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_162_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05337__I _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08855_ _01704_ _03191_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__05709__A1 _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07806_ _02947_ _03058_ _03054_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08648__I _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08786_ _03891_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06382__A1 _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05998_ _01534_ _01541_ _01446_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input13_I i_la_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07737_ _02160_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08659__B1 _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05980__I1 stack\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06168__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07668_ _02952_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ _04369_ _04379_ _04381_ _04382_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06619_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07599_ _02896_ _02889_ _02899_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ _04283_ mem.dff_data_out\[4\] _04318_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ _01171_ _04253_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_139_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05956__B _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07937__A2 _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06631__I _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11162_ _00754_ clknet_leaf_5_clock stack\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__A1 stack\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__I _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _04976_ _04977_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06070__B1 _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11093_ _00685_ clknet_leaf_14_clock net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05247__I _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09942__I _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10044_ _04911_ _04912_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_212_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10427__CLK clknet_leaf_60_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05971__I1 stack\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08114__A2 _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06078__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10946_ _00538_ clknet_leaf_180_clock stack\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05911__S _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07873__A1 _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10877_ _00469_ clknet_leaf_144_clock stack\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09075__B1 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06428__A2 _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06027__B _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09378__A1 _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09338__B _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06541__I _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06970_ _02164_ _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I i_la_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05921_ stack\[8\]\[3\] stack\[9\]\[3\] _01427_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08640_ _03741_ _03637_ _03777_ _03234_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_05852_ _01278_ _01389_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06364__A1 _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10160__A2 _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _01859_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05783_ _01261_ stack\[30\]\[0\] _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08105__A2 _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07522_ mem.mem_dff.code_mem\[26\]\[7\] _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05821__S _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07453_ _02782_ _02775_ _02785_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__I _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06404_ _01935_ _01940_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07384_ _02648_ _02731_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05620__I _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08136__C _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09123_ _04071_ _04146_ _04142_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07616__A1 _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10238__I _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06335_ _01803_ _01806_ _01844_ _01834_ _01838_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06419__A2 _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ _03870_ _04087_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08931__I _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06266_ _01803_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_194_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ _03215_ _03209_ _03205_ stack\[28\]\[1\] _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05217_ _00771_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _01738_ _01739_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08041__A1 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06052__B1 _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__A2 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09956_ _02004_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08907_ _03961_ _03969_ _03983_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09887_ _03261_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08344__A2 _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08838_ _03929_ _03931_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08769_ _03721_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10800_ _00392_ clknet_leaf_163_clock stack\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06107__A1 _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10731_ _00323_ clknet_leaf_50_clock mem.mem_dff.data_mem\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10662_ _00254_ clknet_leaf_78_clock mem.mem_dff.code_mem\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08804__B1 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10593_ _00185_ clknet_leaf_87_clock mem.mem_dff.code_mem\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08280__A1 _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07457__I _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11145_ _00737_ clknet_4_1_0_clock stack\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ _00668_ clknet_leaf_132_clock delay_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10027_ _04885_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06346__A1 _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10929_ _00521_ clknet_leaf_180_clock stack\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06120_ net38 net7 _01654_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06121__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06282__B1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06051_ _01036_ _01033_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_173_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _01891_ _04739_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__A2 _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ _04695_ _04696_ _04697_ _04698_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06953_ _02149_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09515__C _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10118__C1 _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10742__CLK clknet_leaf_163_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _01379_ _01397_ _01425_ _01447_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09672_ _04606_ _04631_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06884_ _02337_ _02334_ _02338_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08623_ _03761_ _03764_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05835_ _01368_ _01378_ _00852_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _03633_ _03707_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05766_ _01264_ stack\[26\]\[2\] _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10892__CLK clknet_leaf_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05560__A2 stack\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ mem.mem_dff.code_mem\[26\]\[3\] _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ _03652_ _03642_ _03648_ stack\[19\]\[2\] _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05697_ _01223_ _01213_ _01208_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07436_ _02742_ _02765_ _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09039__B1 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05312__A2 _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07367_ _02717_ _02718_ _02713_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05863__A3 _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input80_I rambus_wb_dat_i[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__B _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _03847_ _03964_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06318_ stack\[2\]\[3\] _01830_ _01857_ _01759_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08661__I _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ _02662_ _02663_ _02665_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08262__B2 mem.mem_dff.code_mem\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09037_ _04061_ _04067_ _04081_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06249_ _01720_ _01769_ _01790_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A1 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06576__A1 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _04563_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05953__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09514__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06328__A1 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__A2 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05525__I _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07740__I _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05839__B1 _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _00306_ clknet_leaf_30_clock mem.mem_dff.data_mem\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ _00237_ clknet_4_12_0_clock mem.mem_dff.code_mem\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10615__CLK clknet_leaf_106_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08571__I _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10576_ _00168_ clknet_leaf_90_clock mem.mem_dff.code_mem\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08253__B2 mem.mem_dff.data_mem\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06091__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__A1 _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08005__B2 stack\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10765__CLK clknet_leaf_37_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__A1 _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10363__A2 _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11128_ _00720_ clknet_leaf_169_clock stack\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09505__A1 _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07136__B _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _00651_ clknet_leaf_23_clock delay_cycles\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06319__A1 _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10115__A2 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08859__A3 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05620_ _01167_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07650__I _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05542__A2 stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05551_ _01092_ _01095_ _01099_ _01053_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08270_ mem.mem_dff.code_mem\[1\]\[4\] _03355_ _03358_ mem.mem_dff.code_mem\[17\]\[4\]
+ _03356_ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05482_ stack\[23\]\[5\] stack\[20\]\[5\] stack\[21\]\[5\] stack\[22\]\[5\] _01030_
+ _01031_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08492__A1 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08492__B2 stack\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07221_ _02589_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_182_clock clknet_4_4_0_clock clknet_leaf_182_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_220_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08244__A1 mem.mem_dff.code_mem\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _02548_ _02549_ _02551_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08244__B2 mem.mem_dff.code_mem\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06103_ _01632_ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_161_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08795__A2 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__A1 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07083_ _02407_ _02486_ _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06034_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10354__A2 _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__I mem.mem_dff.data_mem\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_120_clock clknet_4_12_0_clock clknet_leaf_120_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07985_ _01587_ _03196_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09724_ _04251_ _04659_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06936_ mem.mem_dff.code_mem\[11\]\[0\] _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10106__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09655_ _04612_ _04613_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06867_ mem.mem_dff.code_mem\[9\]\[1\] _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05908__I1 stack\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_135_clock clknet_4_6_0_clock clknet_leaf_135_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08606_ stack\[3\]\[1\] _03746_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05818_ stack\[16\]\[7\] stack\[17\]\[7\] _01013_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09586_ _04544_ _04545_ _04533_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06730__A1 _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ _02269_ _02261_ _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11070__CLK clknet_leaf_69_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ _03232_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05749_ _01282_ _01287_ _01292_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10638__CLK clknet_leaf_103_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06176__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08483__A1 _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _01689_ _01693_ _01698_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05297__A1 _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07419_ _02531_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10290__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08399_ net122 _02108_ _03578_ _03579_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10430_ _00022_ clknet_leaf_75_clock mem.mem_dff.code_mem\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08391__I _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07038__A2 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10788__CLK clknet_leaf_3_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09983__A1 _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10361_ _01857_ _05154_ _05161_ stack\[17\]\[3\] _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05844__I0 stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ _05111_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10345__A2 _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05221__A1 _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__I _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08710__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08566__I _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07470__I _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07277__A2 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08474__A1 _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10281__A1 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__C _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_146_clock_I clknet_4_5_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10281__B2 stack\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09397__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10628_ _00220_ clknet_leaf_102_clock mem.mem_dff.code_mem\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06814__I _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__A2 _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10033__B2 _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A2 _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10559_ _00151_ clknet_leaf_96_clock mem.mem_dff.code_mem\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A4 _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10336__A2 _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__A2 _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06004__A3 _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07770_ _03030_ _03031_ _03033_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06960__A1 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06721_ _02194_ _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11093__CLK clknet_leaf_14_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04412_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06652_ _02117_ _02155_ _02151_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06712__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05603_ _01144_ stack\[16\]\[7\] stack\[17\]\[7\] _01150_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09371_ net93 _03042_ _03014_ net84 _04281_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06583_ _02018_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_67_clock clknet_4_14_0_clock clknet_leaf_67_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _03512_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05534_ _01012_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__A1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ mem.mem_dff.data_mem\[4\]\[3\] _03101_ _03131_ mem.mem_dff.data_mem\[5\]\[3\]
+ _03381_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__B2 stack\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05465_ _01012_ stack\[28\]\[4\] stack\[29\]\[4\] _01015_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _02589_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__A1 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08184_ _03320_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05396_ _00938_ _00939_ _00947_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07135_ _02537_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05826__I0 stack\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07066_ _02480_ _02471_ _02482_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput230 net230 rambus_wb_sel_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05451__A1 _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06017_ stack\[6\]\[1\] stack\[7\]\[1\] _01374_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10327__A2 _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I i_wb_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09193__A2 _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08940__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ mem.mem_dff.data_mem\[7\]\[6\] _03179_ _03176_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06919_ _02348_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09707_ _04478_ _04666_ _04649_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_210_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07899_ _03073_ _03134_ _03127_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08153__B1 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__CLK clknet_leaf_85_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08386__I _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _04584_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06703__A1 _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05506__A2 stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05357__I2 stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08319__C _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ cycles_per_ms\[15\] _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10263__A1 _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _00005_ clknet_leaf_170_clock stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05690__A1 _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05817__I0 stack\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _05066_ _05148_ _05149_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09708__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10275_ _05057_ _05098_ _05100_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__A2 _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07195__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_clock_I clknet_4_15_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05914__S _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06809__I _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08695__A1 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08695__B2 stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10953__CLK clknet_leaf_149_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10254__B2 stack\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06544__I mem.mem_dff.code_mem\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05250_ net138 _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_128_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05681__A1 _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__A4 _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08940_ _03957_ _04003_ _04010_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10309__A2 _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05984__A2 _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08871_ _03839_ _03947_ _03955_ stack\[26\]\[3\] _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07822_ _03071_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10483__CLK clknet_leaf_56_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07753_ _03019_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06704_ _02193_ _02186_ _02196_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07684_ _02936_ _02960_ _02953_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08686__A1 _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09883__B1 _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05623__I _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09423_ _01827_ _04380_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06635_ mem.mem_dff.code_mem\[3\]\[1\] _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06161__A2 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09354_ _04298_ _01896_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06566_ _02051_ _02085_ _02081_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08438__A1 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__I _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ mem.mem_dff.code_mem\[17\]\[5\] _02562_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10245__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10245__B2 stack\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08989__A2 _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05517_ stack\[11\]\[5\] stack\[8\]\[5\] stack\[9\]\[5\] stack\[10\]\[5\] _01029_
+ _00969_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09285_ mem.sram_enable _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07110__A1 _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06497_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08236_ _02320_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05448_ _00994_ _00996_ _00998_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06454__I _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08167_ mem.mem_dff.code_mem\[8\]\[1\] _02292_ _02700_ mem.mem_dff.code_mem\[22\]\[1\]
+ mem.mem_dff.code_mem\[31\]\[1\] _02957_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_181_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05379_ _00786_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _02523_ _02517_ _02513_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08098_ mem.mem_dff.code_mem\[8\]\[0\] _03292_ _03293_ mem.mem_dff.code_mem\[22\]\[0\]
+ mem.mem_dff.code_mem\[31\]\[0\] _02957_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_107_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__D _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07049_ _02468_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10826__CLK clknet_leaf_169_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09166__A2 _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10060_ _04927_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08913__A2 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__CLK clknet_leaf_42_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06629__I _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10962_ _00554_ clknet_leaf_179_clock stack\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09005__I _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _00485_ clknet_leaf_146_clock stack\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08429__A1 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05415__A1 stack\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10327_ _04191_ _05137_ _05138_ _04915_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A2 _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10258_ _03908_ _05086_ _05071_ _03733_ _05087_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08904__A2 _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ _04950_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05274__S0 _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06539__I _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__A1 _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08668__B2 stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06983__B _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06420_ net14 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11131__CLK clknet_leaf_173_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07891__A2 _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10227__A1 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06351_ _01861_ _01641_ _01889_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09093__A1 _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__B2 stack\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05302_ _00855_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09070_ _03228_ _04085_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06282_ _01720_ _01800_ _01819_ _01822_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08840__A1 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__B2 stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08021_ _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05233_ _00783_ _00787_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10849__CLK clknet_leaf_162_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05406__A1 _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05257__I1 stack\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _04857_ _04860_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05957__A2 stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09148__A2 _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08923_ _03996_ _03991_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10999__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08854_ _01928_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_85_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05709__A2 _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07805_ mem.mem_dff.data_mem\[2\]\[5\] _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _01639_ _03807_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05997_ _01380_ _01537_ _01540_ _01436_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07736_ _03005_ _03002_ _03006_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07054__B _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08659__A1 _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09856__B1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08659__B2 stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ _02840_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__A1 _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06618_ _01997_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09406_ _04323_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ _02870_ _02890_ _02898_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05893__A1 _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06549_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09337_ _04316_ _04317_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09084__A1 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_clock_I clknet_4_8_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09268_ net77 net193 mem.dff_data_ready mem.io_data_ready _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07634__A2 _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08831__A1 stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output197_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08219_ mem.mem_dff.data_mem\[2\]\[2\] _03044_ _03375_ mem.mem_dff.data_mem\[6\]\[2\]
+ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_154_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09199_ _04180_ _04195_ _04202_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06912__I _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09428__C _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _00753_ clknet_leaf_166_clock stack\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05528__I _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10112_ _04587_ _04963_ _04943_ _01255_ net153 _04939_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05799__I2 stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__A2 _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11092_ _00684_ clknet_leaf_14_clock net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11004__CLK clknet_leaf_129_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10043_ delay_counter\[7\] _04674_ _04899_ _01169_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08898__A1 _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11154__CLK clknet_leaf_191_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10945_ _00537_ clknet_leaf_149_clock stack\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07322__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _00468_ clknet_leaf_192_clock stack\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09075__A1 _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09075__B2 stack\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09378__A2 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07139__B _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06061__A1 _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ stack\[10\]\[3\] stack\[11\]\[3\] _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08889__A1 _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05851_ _01390_ _01392_ _01393_ _01394_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_212_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11175__I clknet_opt_4_1_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08570_ stack\[31\]\[4\] _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05782_ stack\[31\]\[0\] _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07521_ _02837_ _02830_ _02838_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10521__CLK clknet_leaf_112_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__A1 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02755_ _02776_ _02784_ _02785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06403_ _01937_ _01938_ _01939_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_204_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ _04146_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10671__CLK clknet_leaf_59_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06334_ _01834_ _01844_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08813__A1 stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05627__A1 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _04091_ _04094_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06265_ _01579_ _01805_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07828__I mem.mem_dff.data_mem\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08004_ _03214_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05216_ _00767_ _00770_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06196_ _00839_ _01578_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11027__CLK clknet_leaf_17_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05348__I _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ _04840_ _04849_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _03844_ _03971_ _03979_ stack\[10\]\[5\] _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09886_ _04791_ _04797_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _03224_ _03913_ _03930_ net148 _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _03877_ _03878_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output112_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _02143_ _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_199_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _01587_ _03196_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10730_ _00322_ clknet_leaf_64_clock mem.mem_dff.data_mem\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08394__I _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08327__C _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _00253_ clknet_leaf_57_clock mem.mem_dff.code_mem\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09057__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10592_ _00184_ clknet_leaf_87_clock mem.mem_dff.code_mem\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08804__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__B2 stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05618__A1 _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08280__A2 _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11144_ _00736_ clknet_leaf_177_clock stack\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07791__A1 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11075_ _00667_ clknet_4_9_0_clock delay_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07473__I mem.mem_dff.code_mem\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10026_ _04894_ _04895_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10544__CLK clknet_leaf_97_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06089__I _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09296__A1 _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10694__CLK clknet_4_14_0_clock vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06817__I mem.mem_dff.code_mem\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10928_ _00520_ clknet_leaf_147_clock stack\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10859_ _00451_ clknet_leaf_0_clock stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05609__A1 _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06050_ _01581_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05468__S0 _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06952_ mem.mem_dff.code_mem\[11\]\[3\] _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09740_ cycles_per_ms\[7\] _04577_ _04592_ _04593_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

