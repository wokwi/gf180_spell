* NGSPICE file created from user_project_wrapper.ext - technology: gf180mcuC

* Black-box entry subcircuit for rambus abstract view
.subckt rambus rambus_wb_ack_o rambus_wb_addr_i[0] rambus_wb_addr_i[1] rambus_wb_addr_i[2]
+ rambus_wb_addr_i[3] rambus_wb_addr_i[4] rambus_wb_addr_i[5] rambus_wb_addr_i[6]
+ rambus_wb_addr_i[7] rambus_wb_addr_i[8] rambus_wb_clk_i rambus_wb_cyc_i rambus_wb_dat_i[0]
+ rambus_wb_dat_i[10] rambus_wb_dat_i[11] rambus_wb_dat_i[12] rambus_wb_dat_i[13]
+ rambus_wb_dat_i[14] rambus_wb_dat_i[15] rambus_wb_dat_i[16] rambus_wb_dat_i[17]
+ rambus_wb_dat_i[18] rambus_wb_dat_i[19] rambus_wb_dat_i[1] rambus_wb_dat_i[20] rambus_wb_dat_i[21]
+ rambus_wb_dat_i[22] rambus_wb_dat_i[23] rambus_wb_dat_i[24] rambus_wb_dat_i[25]
+ rambus_wb_dat_i[26] rambus_wb_dat_i[27] rambus_wb_dat_i[28] rambus_wb_dat_i[29]
+ rambus_wb_dat_i[2] rambus_wb_dat_i[30] rambus_wb_dat_i[31] rambus_wb_dat_i[3] rambus_wb_dat_i[4]
+ rambus_wb_dat_i[5] rambus_wb_dat_i[6] rambus_wb_dat_i[7] rambus_wb_dat_i[8] rambus_wb_dat_i[9]
+ rambus_wb_dat_o[0] rambus_wb_dat_o[10] rambus_wb_dat_o[11] rambus_wb_dat_o[12] rambus_wb_dat_o[13]
+ rambus_wb_dat_o[14] rambus_wb_dat_o[15] rambus_wb_dat_o[16] rambus_wb_dat_o[17]
+ rambus_wb_dat_o[18] rambus_wb_dat_o[19] rambus_wb_dat_o[1] rambus_wb_dat_o[20] rambus_wb_dat_o[21]
+ rambus_wb_dat_o[22] rambus_wb_dat_o[23] rambus_wb_dat_o[24] rambus_wb_dat_o[25]
+ rambus_wb_dat_o[26] rambus_wb_dat_o[27] rambus_wb_dat_o[28] rambus_wb_dat_o[29]
+ rambus_wb_dat_o[2] rambus_wb_dat_o[30] rambus_wb_dat_o[31] rambus_wb_dat_o[3] rambus_wb_dat_o[4]
+ rambus_wb_dat_o[5] rambus_wb_dat_o[6] rambus_wb_dat_o[7] rambus_wb_dat_o[8] rambus_wb_dat_o[9]
+ rambus_wb_rst_i rambus_wb_sel_i[0] rambus_wb_sel_i[1] rambus_wb_sel_i[2] rambus_wb_sel_i[3]
+ rambus_wb_stb_i rambus_wb_we_i vdd vss
.ends

* Black-box entry subcircuit for spell abstract view
.subckt spell clock i_la_addr[0] i_la_addr[1] i_la_addr[2] i_la_addr[3] i_la_addr[4]
+ i_la_addr[5] i_la_addr[6] i_la_data[0] i_la_data[1] i_la_data[2] i_la_data[3] i_la_data[4]
+ i_la_data[5] i_la_data[6] i_la_data[7] i_la_wb_disable i_la_write i_wb_addr[0] i_wb_addr[10]
+ i_wb_addr[11] i_wb_addr[12] i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16]
+ i_wb_addr[17] i_wb_addr[18] i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21]
+ i_wb_addr[22] i_wb_addr[23] i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27]
+ i_wb_addr[28] i_wb_addr[29] i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3]
+ i_wb_addr[4] i_wb_addr[5] i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc
+ i_wb_data[0] i_wb_data[10] i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14]
+ i_wb_data[15] i_wb_data[16] i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1]
+ i_wb_data[20] i_wb_data[21] i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25]
+ i_wb_data[26] i_wb_data[27] i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30]
+ i_wb_data[31] i_wb_data[3] i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8]
+ i_wb_data[9] i_wb_stb i_wb_we interrupt io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_oeb[0] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3]
+ la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ o_wb_ack o_wb_data[0] o_wb_data[10] o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14]
+ o_wb_data[15] o_wb_data[16] o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1]
+ o_wb_data[20] o_wb_data[21] o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25]
+ o_wb_data[26] o_wb_data[27] o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30]
+ o_wb_data[31] o_wb_data[3] o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8]
+ o_wb_data[9] rambus_wb_ack_i rambus_wb_addr_o[0] rambus_wb_addr_o[1] rambus_wb_addr_o[2]
+ rambus_wb_addr_o[3] rambus_wb_addr_o[4] rambus_wb_addr_o[5] rambus_wb_addr_o[6]
+ rambus_wb_addr_o[7] rambus_wb_addr_o[8] rambus_wb_addr_o[9] rambus_wb_clk_o rambus_wb_cyc_o
+ rambus_wb_dat_i[0] rambus_wb_dat_i[10] rambus_wb_dat_i[11] rambus_wb_dat_i[12] rambus_wb_dat_i[13]
+ rambus_wb_dat_i[14] rambus_wb_dat_i[15] rambus_wb_dat_i[16] rambus_wb_dat_i[17]
+ rambus_wb_dat_i[18] rambus_wb_dat_i[19] rambus_wb_dat_i[1] rambus_wb_dat_i[20] rambus_wb_dat_i[21]
+ rambus_wb_dat_i[22] rambus_wb_dat_i[23] rambus_wb_dat_i[24] rambus_wb_dat_i[25]
+ rambus_wb_dat_i[26] rambus_wb_dat_i[27] rambus_wb_dat_i[28] rambus_wb_dat_i[29]
+ rambus_wb_dat_i[2] rambus_wb_dat_i[30] rambus_wb_dat_i[31] rambus_wb_dat_i[3] rambus_wb_dat_i[4]
+ rambus_wb_dat_i[5] rambus_wb_dat_i[6] rambus_wb_dat_i[7] rambus_wb_dat_i[8] rambus_wb_dat_i[9]
+ rambus_wb_dat_o[0] rambus_wb_dat_o[10] rambus_wb_dat_o[11] rambus_wb_dat_o[12] rambus_wb_dat_o[13]
+ rambus_wb_dat_o[14] rambus_wb_dat_o[15] rambus_wb_dat_o[16] rambus_wb_dat_o[17]
+ rambus_wb_dat_o[18] rambus_wb_dat_o[19] rambus_wb_dat_o[1] rambus_wb_dat_o[20] rambus_wb_dat_o[21]
+ rambus_wb_dat_o[22] rambus_wb_dat_o[23] rambus_wb_dat_o[24] rambus_wb_dat_o[25]
+ rambus_wb_dat_o[26] rambus_wb_dat_o[27] rambus_wb_dat_o[28] rambus_wb_dat_o[29]
+ rambus_wb_dat_o[2] rambus_wb_dat_o[30] rambus_wb_dat_o[31] rambus_wb_dat_o[3] rambus_wb_dat_o[4]
+ rambus_wb_dat_o[5] rambus_wb_dat_o[6] rambus_wb_dat_o[7] rambus_wb_dat_o[8] rambus_wb_dat_o[9]
+ rambus_wb_rst_o rambus_wb_sel_o[0] rambus_wb_sel_o[1] rambus_wb_sel_o[2] rambus_wb_sel_o[3]
+ rambus_wb_stb_o rambus_wb_we_o reset vdd vss
.ends

.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xrambus0 rambus_wb_ack rambus_wb_addr\[0\] rambus_wb_addr\[1\] rambus_wb_addr\[2\]
+ rambus_wb_addr\[3\] rambus_wb_addr\[4\] rambus_wb_addr\[5\] rambus_wb_addr\[6\]
+ rambus_wb_addr\[7\] rambus_wb_addr\[8\] rambus_wb_clk rambus_wb_cyc rambus_wb_dat_i\[0\]
+ rambus_wb_dat_i\[10\] rambus_wb_dat_i\[11\] rambus_wb_dat_i\[12\] rambus_wb_dat_i\[13\]
+ rambus_wb_dat_i\[14\] rambus_wb_dat_i\[15\] rambus_wb_dat_i\[16\] rambus_wb_dat_i\[17\]
+ rambus_wb_dat_i\[18\] rambus_wb_dat_i\[19\] rambus_wb_dat_i\[1\] rambus_wb_dat_i\[20\]
+ rambus_wb_dat_i\[21\] rambus_wb_dat_i\[22\] rambus_wb_dat_i\[23\] rambus_wb_dat_i\[24\]
+ rambus_wb_dat_i\[25\] rambus_wb_dat_i\[26\] rambus_wb_dat_i\[27\] rambus_wb_dat_i\[28\]
+ rambus_wb_dat_i\[29\] rambus_wb_dat_i\[2\] rambus_wb_dat_i\[30\] rambus_wb_dat_i\[31\]
+ rambus_wb_dat_i\[3\] rambus_wb_dat_i\[4\] rambus_wb_dat_i\[5\] rambus_wb_dat_i\[6\]
+ rambus_wb_dat_i\[7\] rambus_wb_dat_i\[8\] rambus_wb_dat_i\[9\] rambus_wb_dat_o\[0\]
+ rambus_wb_dat_o\[10\] rambus_wb_dat_o\[11\] rambus_wb_dat_o\[12\] rambus_wb_dat_o\[13\]
+ rambus_wb_dat_o\[14\] rambus_wb_dat_o\[15\] rambus_wb_dat_o\[16\] rambus_wb_dat_o\[17\]
+ rambus_wb_dat_o\[18\] rambus_wb_dat_o\[19\] rambus_wb_dat_o\[1\] rambus_wb_dat_o\[20\]
+ rambus_wb_dat_o\[21\] rambus_wb_dat_o\[22\] rambus_wb_dat_o\[23\] rambus_wb_dat_o\[24\]
+ rambus_wb_dat_o\[25\] rambus_wb_dat_o\[26\] rambus_wb_dat_o\[27\] rambus_wb_dat_o\[28\]
+ rambus_wb_dat_o\[29\] rambus_wb_dat_o\[2\] rambus_wb_dat_o\[30\] rambus_wb_dat_o\[31\]
+ rambus_wb_dat_o\[3\] rambus_wb_dat_o\[4\] rambus_wb_dat_o\[5\] rambus_wb_dat_o\[6\]
+ rambus_wb_dat_o\[7\] rambus_wb_dat_o\[8\] rambus_wb_dat_o\[9\] rambus_wb_rst rambus_wb_sel\[0\]
+ rambus_wb_sel\[1\] rambus_wb_sel\[2\] rambus_wb_sel\[3\] rambus_wb_stb rambus_wb_we
+ vdd vss rambus
Xspell wb_clk_i la_data_in[8] la_data_in[9] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[1] la_data_in[2]
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_stb_i wbs_we_i user_irq[0] io_in[8] io_in[9]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_oeb[8] io_oeb[9]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_out[8] io_out[9]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] la_data_out[0]
+ la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[3] la_data_out[4] la_data_out[5]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] wbs_ack_o wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ rambus_wb_ack rambus_wb_addr\[0\] rambus_wb_addr\[1\] rambus_wb_addr\[2\] rambus_wb_addr\[3\]
+ rambus_wb_addr\[4\] rambus_wb_addr\[5\] rambus_wb_addr\[6\] rambus_wb_addr\[7\]
+ rambus_wb_addr\[8\] spell/rambus_wb_addr_o[9] rambus_wb_clk rambus_wb_cyc rambus_wb_dat_o\[0\]
+ rambus_wb_dat_o\[10\] rambus_wb_dat_o\[11\] rambus_wb_dat_o\[12\] rambus_wb_dat_o\[13\]
+ rambus_wb_dat_o\[14\] rambus_wb_dat_o\[15\] rambus_wb_dat_o\[16\] rambus_wb_dat_o\[17\]
+ rambus_wb_dat_o\[18\] rambus_wb_dat_o\[19\] rambus_wb_dat_o\[1\] rambus_wb_dat_o\[20\]
+ rambus_wb_dat_o\[21\] rambus_wb_dat_o\[22\] rambus_wb_dat_o\[23\] rambus_wb_dat_o\[24\]
+ rambus_wb_dat_o\[25\] rambus_wb_dat_o\[26\] rambus_wb_dat_o\[27\] rambus_wb_dat_o\[28\]
+ rambus_wb_dat_o\[29\] rambus_wb_dat_o\[2\] rambus_wb_dat_o\[30\] rambus_wb_dat_o\[31\]
+ rambus_wb_dat_o\[3\] rambus_wb_dat_o\[4\] rambus_wb_dat_o\[5\] rambus_wb_dat_o\[6\]
+ rambus_wb_dat_o\[7\] rambus_wb_dat_o\[8\] rambus_wb_dat_o\[9\] rambus_wb_dat_i\[0\]
+ rambus_wb_dat_i\[10\] rambus_wb_dat_i\[11\] rambus_wb_dat_i\[12\] rambus_wb_dat_i\[13\]
+ rambus_wb_dat_i\[14\] rambus_wb_dat_i\[15\] rambus_wb_dat_i\[16\] rambus_wb_dat_i\[17\]
+ rambus_wb_dat_i\[18\] rambus_wb_dat_i\[19\] rambus_wb_dat_i\[1\] rambus_wb_dat_i\[20\]
+ rambus_wb_dat_i\[21\] rambus_wb_dat_i\[22\] rambus_wb_dat_i\[23\] rambus_wb_dat_i\[24\]
+ rambus_wb_dat_i\[25\] rambus_wb_dat_i\[26\] rambus_wb_dat_i\[27\] rambus_wb_dat_i\[28\]
+ rambus_wb_dat_i\[29\] rambus_wb_dat_i\[2\] rambus_wb_dat_i\[30\] rambus_wb_dat_i\[31\]
+ rambus_wb_dat_i\[3\] rambus_wb_dat_i\[4\] rambus_wb_dat_i\[5\] rambus_wb_dat_i\[6\]
+ rambus_wb_dat_i\[7\] rambus_wb_dat_i\[8\] rambus_wb_dat_i\[9\] rambus_wb_rst rambus_wb_sel\[0\]
+ rambus_wb_sel\[1\] rambus_wb_sel\[2\] rambus_wb_sel\[3\] rambus_wb_stb rambus_wb_we
+ wb_rst_i vdd vss spell
.ends

